module testbench();

    // Input signals
    logic        clk;
    logic [63:0] word;
    logic        pe;
    logic        tkk;

    // Output signals
    logic  [3:0] ir;
    logic  [7:0] op;
    logic        extop;
    logic [19:0] addr;

    // Device under test
    standardizer dut(clk, word, pe, tkk,
        ir, op, extop, addr);

    // Status
    bit fail;

initial begin
$display("------------------------");
$dumpfile("test.vcd");
$dumpvars();
fail = 0;
clk = 0;

// ***************************************************
// * Test vectors for micro-BESM instruction decoder *
// ***************************************************
// 0000000000000001:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 0: ir 'h%h !== 'h0", ir); end	// Vector No: 0
assert (op === 'h00) else begin fail = 1; $display("Error 1: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000001:0:1:0:00:0:00001:
//------------------------

#2;
word <= 'h0000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 2
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4: ir 'h%h !== 'h0", ir); end	// Vector No: 1
assert (op === 'h00) else begin fail = 1; $display("Error 5: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 7: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000000000001:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 3
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 8: ir 'h%h !== 'h0", ir); end	// Vector No: 2
assert (op === 'h00) else begin fail = 1; $display("Error 9: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 10: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 11: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000001:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 4
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 12: ir 'h%h !== 'h0", ir); end	// Vector No: 3
assert (op === 'h00) else begin fail = 1; $display("Error 13: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 14: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 15: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000002:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000002;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 5
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 16: ir 'h%h !== 'h0", ir); end	// Vector No: 4
assert (op === 'h00) else begin fail = 1; $display("Error 17: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 18: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 19: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000002:0:1:0:00:0:00002:
//------------------------

#2;
word <= 'h0000000000000002;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 6
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 20: ir 'h%h !== 'h0", ir); end	// Vector No: 5
assert (op === 'h00) else begin fail = 1; $display("Error 21: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 22: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 23: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000000000002:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000002;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 7
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 24: ir 'h%h !== 'h0", ir); end	// Vector No: 6
assert (op === 'h00) else begin fail = 1; $display("Error 25: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 26: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 27: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000002:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000002;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 8
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 28: ir 'h%h !== 'h0", ir); end	// Vector No: 7
assert (op === 'h00) else begin fail = 1; $display("Error 29: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 30: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 31: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000004:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000004;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 9
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 32: ir 'h%h !== 'h0", ir); end	// Vector No: 8
assert (op === 'h00) else begin fail = 1; $display("Error 33: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 34: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 35: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000004:0:1:0:00:0:00004:
//------------------------

#2;
word <= 'h0000000000000004;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 10
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 36: ir 'h%h !== 'h0", ir); end	// Vector No: 9
assert (op === 'h00) else begin fail = 1; $display("Error 37: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 38: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 39: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000000000004:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000004;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 11
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 40: ir 'h%h !== 'h0", ir); end	// Vector No: 10
assert (op === 'h00) else begin fail = 1; $display("Error 41: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 42: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 43: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000004:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000004;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 12
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 44: ir 'h%h !== 'h0", ir); end	// Vector No: 11
assert (op === 'h00) else begin fail = 1; $display("Error 45: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 46: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 47: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000008:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000008;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 13
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 48: ir 'h%h !== 'h0", ir); end	// Vector No: 12
assert (op === 'h00) else begin fail = 1; $display("Error 49: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 50: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 51: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000008:0:1:0:00:0:00008:
//------------------------

#2;
word <= 'h0000000000000008;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 14
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 52: ir 'h%h !== 'h0", ir); end	// Vector No: 13
assert (op === 'h00) else begin fail = 1; $display("Error 53: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 54: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 55: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000000000008:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000008;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 15
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 56: ir 'h%h !== 'h0", ir); end	// Vector No: 14
assert (op === 'h00) else begin fail = 1; $display("Error 57: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 58: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 59: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000008:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000008;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 16
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 60: ir 'h%h !== 'h0", ir); end	// Vector No: 15
assert (op === 'h00) else begin fail = 1; $display("Error 61: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 62: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 63: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000010:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 17
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 64: ir 'h%h !== 'h0", ir); end	// Vector No: 16
assert (op === 'h00) else begin fail = 1; $display("Error 65: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 66: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 67: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000010:0:1:0:00:0:00010:
//------------------------

#2;
word <= 'h0000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 18
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 68: ir 'h%h !== 'h0", ir); end	// Vector No: 17
assert (op === 'h00) else begin fail = 1; $display("Error 69: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 70: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 71: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000000000010:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 19
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 72: ir 'h%h !== 'h0", ir); end	// Vector No: 18
assert (op === 'h00) else begin fail = 1; $display("Error 73: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 74: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 75: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000010:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 20
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 76: ir 'h%h !== 'h0", ir); end	// Vector No: 19
assert (op === 'h00) else begin fail = 1; $display("Error 77: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 78: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 79: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000020:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000020;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 21
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 80: ir 'h%h !== 'h0", ir); end	// Vector No: 20
assert (op === 'h00) else begin fail = 1; $display("Error 81: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 82: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 83: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000020:0:1:0:00:0:00020:
//------------------------

#2;
word <= 'h0000000000000020;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 22
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 84: ir 'h%h !== 'h0", ir); end	// Vector No: 21
assert (op === 'h00) else begin fail = 1; $display("Error 85: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 86: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 87: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000000000020:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000020;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 23
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 88: ir 'h%h !== 'h0", ir); end	// Vector No: 22
assert (op === 'h00) else begin fail = 1; $display("Error 89: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 90: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 91: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000020:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000020;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 24
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 92: ir 'h%h !== 'h0", ir); end	// Vector No: 23
assert (op === 'h00) else begin fail = 1; $display("Error 93: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 94: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 95: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000040:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000040;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 25
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 96: ir 'h%h !== 'h0", ir); end	// Vector No: 24
assert (op === 'h00) else begin fail = 1; $display("Error 97: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 98: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 99: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000040:0:1:0:00:0:00040:
//------------------------

#2;
word <= 'h0000000000000040;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 26
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 100: ir 'h%h !== 'h0", ir); end	// Vector No: 25
assert (op === 'h00) else begin fail = 1; $display("Error 101: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 102: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 103: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000000000040:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000040;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 27
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 104: ir 'h%h !== 'h0", ir); end	// Vector No: 26
assert (op === 'h00) else begin fail = 1; $display("Error 105: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 106: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 107: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000040:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000040;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 28
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 108: ir 'h%h !== 'h0", ir); end	// Vector No: 27
assert (op === 'h00) else begin fail = 1; $display("Error 109: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 110: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 111: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000080:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000080;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 29
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 112: ir 'h%h !== 'h0", ir); end	// Vector No: 28
assert (op === 'h00) else begin fail = 1; $display("Error 113: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 114: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 115: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000080:0:1:0:00:0:00080:
//------------------------

#2;
word <= 'h0000000000000080;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 30
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 116: ir 'h%h !== 'h0", ir); end	// Vector No: 29
assert (op === 'h00) else begin fail = 1; $display("Error 117: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 118: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 119: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000000000080:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000080;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 31
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 120: ir 'h%h !== 'h0", ir); end	// Vector No: 30
assert (op === 'h00) else begin fail = 1; $display("Error 121: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 122: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 123: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000080:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000080;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 32
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 124: ir 'h%h !== 'h0", ir); end	// Vector No: 31
assert (op === 'h00) else begin fail = 1; $display("Error 125: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 126: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 127: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000100:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 33
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 128: ir 'h%h !== 'h0", ir); end	// Vector No: 32
assert (op === 'h00) else begin fail = 1; $display("Error 129: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 130: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 131: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000100:0:1:0:00:0:00100:
//------------------------

#2;
word <= 'h0000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 34
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 132: ir 'h%h !== 'h0", ir); end	// Vector No: 33
assert (op === 'h00) else begin fail = 1; $display("Error 133: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 134: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 135: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000000000000100:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 35
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 136: ir 'h%h !== 'h0", ir); end	// Vector No: 34
assert (op === 'h00) else begin fail = 1; $display("Error 137: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 138: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 139: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000100:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 36
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 140: ir 'h%h !== 'h0", ir); end	// Vector No: 35
assert (op === 'h00) else begin fail = 1; $display("Error 141: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 142: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 143: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000200:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000200;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 37
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 144: ir 'h%h !== 'h0", ir); end	// Vector No: 36
assert (op === 'h00) else begin fail = 1; $display("Error 145: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 146: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 147: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000200:0:1:0:00:0:00200:
//------------------------

#2;
word <= 'h0000000000000200;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 38
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 148: ir 'h%h !== 'h0", ir); end	// Vector No: 37
assert (op === 'h00) else begin fail = 1; $display("Error 149: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 150: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 151: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000000000000200:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000200;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 39
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 152: ir 'h%h !== 'h0", ir); end	// Vector No: 38
assert (op === 'h00) else begin fail = 1; $display("Error 153: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 154: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 155: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000200:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000200;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 40
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 156: ir 'h%h !== 'h0", ir); end	// Vector No: 39
assert (op === 'h00) else begin fail = 1; $display("Error 157: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 158: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 159: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000400:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000400;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 41
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 160: ir 'h%h !== 'h0", ir); end	// Vector No: 40
assert (op === 'h00) else begin fail = 1; $display("Error 161: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 162: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 163: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000400:0:1:0:00:0:00400:
//------------------------

#2;
word <= 'h0000000000000400;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 42
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 164: ir 'h%h !== 'h0", ir); end	// Vector No: 41
assert (op === 'h00) else begin fail = 1; $display("Error 165: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 166: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 167: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000000000000400:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000400;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 43
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 168: ir 'h%h !== 'h0", ir); end	// Vector No: 42
assert (op === 'h00) else begin fail = 1; $display("Error 169: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 170: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 171: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000400:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000400;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 44
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 172: ir 'h%h !== 'h0", ir); end	// Vector No: 43
assert (op === 'h00) else begin fail = 1; $display("Error 173: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 174: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 175: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000800:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000800;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 45
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 176: ir 'h%h !== 'h0", ir); end	// Vector No: 44
assert (op === 'h00) else begin fail = 1; $display("Error 177: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 178: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 179: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000800:0:1:0:00:0:00800:
//------------------------

#2;
word <= 'h0000000000000800;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 46
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 180: ir 'h%h !== 'h0", ir); end	// Vector No: 45
assert (op === 'h00) else begin fail = 1; $display("Error 181: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 182: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 183: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000000000000800:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000800;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 47
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 184: ir 'h%h !== 'h0", ir); end	// Vector No: 46
assert (op === 'h00) else begin fail = 1; $display("Error 185: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 186: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 187: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000000800:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000000800;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 48
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 188: ir 'h%h !== 'h0", ir); end	// Vector No: 47
assert (op === 'h00) else begin fail = 1; $display("Error 189: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 190: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 191: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000001000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 49
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 192: ir 'h%h !== 'h0", ir); end	// Vector No: 48
assert (op === 'h00) else begin fail = 1; $display("Error 193: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 194: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 195: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000001000:0:1:0:00:0:01000:
//------------------------

#2;
word <= 'h0000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 50
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 196: ir 'h%h !== 'h0", ir); end	// Vector No: 49
assert (op === 'h00) else begin fail = 1; $display("Error 197: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 198: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 199: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000000000001000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 51
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 200: ir 'h%h !== 'h0", ir); end	// Vector No: 50
assert (op === 'h00) else begin fail = 1; $display("Error 201: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 202: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 203: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000001000:1:1:0:00:0:00001:
//------------------------

#2;
word <= 'h0000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 52
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 204: ir 'h%h !== 'h0", ir); end	// Vector No: 51
assert (op === 'h00) else begin fail = 1; $display("Error 205: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 206: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 207: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000000002000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000002000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 53
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 208: ir 'h%h !== 'h0", ir); end	// Vector No: 52
assert (op === 'h00) else begin fail = 1; $display("Error 209: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 210: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 211: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000002000:0:1:0:00:0:02000:
//------------------------

#2;
word <= 'h0000000000002000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 54
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 212: ir 'h%h !== 'h0", ir); end	// Vector No: 53
assert (op === 'h00) else begin fail = 1; $display("Error 213: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 214: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 215: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000000000002000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000002000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 55
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 216: ir 'h%h !== 'h0", ir); end	// Vector No: 54
assert (op === 'h00) else begin fail = 1; $display("Error 217: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 218: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 219: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000002000:1:1:0:00:0:00002:
//------------------------

#2;
word <= 'h0000000000002000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 56
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 220: ir 'h%h !== 'h0", ir); end	// Vector No: 55
assert (op === 'h00) else begin fail = 1; $display("Error 221: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 222: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 223: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000000004000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000004000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 57
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 224: ir 'h%h !== 'h0", ir); end	// Vector No: 56
assert (op === 'h00) else begin fail = 1; $display("Error 225: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 226: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 227: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000004000:0:1:0:00:0:04000:
//------------------------

#2;
word <= 'h0000000000004000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 58
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 228: ir 'h%h !== 'h0", ir); end	// Vector No: 57
assert (op === 'h00) else begin fail = 1; $display("Error 229: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 230: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 231: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000000000004000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000004000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 59
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 232: ir 'h%h !== 'h0", ir); end	// Vector No: 58
assert (op === 'h00) else begin fail = 1; $display("Error 233: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 234: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 235: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000004000:1:1:0:00:0:00004:
//------------------------

#2;
word <= 'h0000000000004000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 60
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 236: ir 'h%h !== 'h0", ir); end	// Vector No: 59
assert (op === 'h00) else begin fail = 1; $display("Error 237: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 238: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 239: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000000008000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000008000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 61
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 240: ir 'h%h !== 'h0", ir); end	// Vector No: 60
assert (op === 'h00) else begin fail = 1; $display("Error 241: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 242: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 243: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000008000:0:1:0:00:0:08000:
//------------------------

#2;
word <= 'h0000000000008000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 62
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 244: ir 'h%h !== 'h0", ir); end	// Vector No: 61
assert (op === 'h00) else begin fail = 1; $display("Error 245: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 246: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 247: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000000000008000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000008000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 63
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 248: ir 'h%h !== 'h0", ir); end	// Vector No: 62
assert (op === 'h00) else begin fail = 1; $display("Error 249: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 250: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 251: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000008000:1:1:0:00:0:00008:
//------------------------

#2;
word <= 'h0000000000008000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 64
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 252: ir 'h%h !== 'h0", ir); end	// Vector No: 63
assert (op === 'h00) else begin fail = 1; $display("Error 253: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 254: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 255: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000000010000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 65
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 256: ir 'h%h !== 'h0", ir); end	// Vector No: 64
assert (op === 'h00) else begin fail = 1; $display("Error 257: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 258: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 259: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000010000:0:1:0:00:0:10000:
//------------------------

#2;
word <= 'h0000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 66
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 260: ir 'h%h !== 'h0", ir); end	// Vector No: 65
assert (op === 'h00) else begin fail = 1; $display("Error 261: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 262: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 263: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0000000000010000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 67
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 264: ir 'h%h !== 'h0", ir); end	// Vector No: 66
assert (op === 'h00) else begin fail = 1; $display("Error 265: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 266: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 267: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000010000:1:1:0:00:0:00010:
//------------------------

#2;
word <= 'h0000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 68
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 268: ir 'h%h !== 'h0", ir); end	// Vector No: 67
assert (op === 'h00) else begin fail = 1; $display("Error 269: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 270: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 271: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000000020000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000020000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 69
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 272: ir 'h%h !== 'h0", ir); end	// Vector No: 68
assert (op === 'h00) else begin fail = 1; $display("Error 273: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 274: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 275: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000020000:0:1:0:00:0:20000:
//------------------------

#2;
word <= 'h0000000000020000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 70
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 276: ir 'h%h !== 'h0", ir); end	// Vector No: 69
assert (op === 'h00) else begin fail = 1; $display("Error 277: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 278: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 279: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0000000000020000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000020000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 71
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 280: ir 'h%h !== 'h0", ir); end	// Vector No: 70
assert (op === 'h00) else begin fail = 1; $display("Error 281: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 282: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 283: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000020000:1:1:0:00:0:00020:
//------------------------

#2;
word <= 'h0000000000020000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 72
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 284: ir 'h%h !== 'h0", ir); end	// Vector No: 71
assert (op === 'h00) else begin fail = 1; $display("Error 285: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 286: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 287: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000000040000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000040000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 73
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 288: ir 'h%h !== 'h0", ir); end	// Vector No: 72
assert (op === 'h00) else begin fail = 1; $display("Error 289: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 290: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 291: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000040000:0:1:0:00:0:40000:
//------------------------

#2;
word <= 'h0000000000040000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 74
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 292: ir 'h%h !== 'h0", ir); end	// Vector No: 73
assert (op === 'h00) else begin fail = 1; $display("Error 293: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 294: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 295: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0000000000040000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000040000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 75
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 296: ir 'h%h !== 'h0", ir); end	// Vector No: 74
assert (op === 'h00) else begin fail = 1; $display("Error 297: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 298: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 299: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000040000:1:1:0:00:0:00040:
//------------------------

#2;
word <= 'h0000000000040000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 76
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 300: ir 'h%h !== 'h0", ir); end	// Vector No: 75
assert (op === 'h00) else begin fail = 1; $display("Error 301: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 302: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 303: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000000080000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000080000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 77
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 304: ir 'h%h !== 'h0", ir); end	// Vector No: 76
assert (op === 'h00) else begin fail = 1; $display("Error 305: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 306: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 307: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000080000:0:1:0:00:0:80000:
//------------------------

#2;
word <= 'h0000000000080000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 78
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 308: ir 'h%h !== 'h0", ir); end	// Vector No: 77
assert (op === 'h00) else begin fail = 1; $display("Error 309: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 310: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 311: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0000000000080000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000080000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 79
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 312: ir 'h%h !== 'h0", ir); end	// Vector No: 78
assert (op === 'h00) else begin fail = 1; $display("Error 313: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 314: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 315: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000080000:1:1:0:00:0:00080:
//------------------------

#2;
word <= 'h0000000000080000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 80
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 316: ir 'h%h !== 'h0", ir); end	// Vector No: 79
assert (op === 'h00) else begin fail = 1; $display("Error 317: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 318: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 319: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000000100000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 81
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 320: ir 'h%h !== 'h0", ir); end	// Vector No: 80
assert (op === 'h00) else begin fail = 1; $display("Error 321: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 322: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 323: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000100000:0:1:0:01:0:00000:
//------------------------

#2;
word <= 'h0000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 82
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 324: ir 'h%h !== 'h0", ir); end	// Vector No: 81
assert (op === 'h01) else begin fail = 1; $display("Error 325: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 326: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 327: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000100000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 83
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 328: ir 'h%h !== 'h0", ir); end	// Vector No: 82
assert (op === 'h00) else begin fail = 1; $display("Error 329: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 330: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 331: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000100000:1:1:0:00:0:00100:
//------------------------

#2;
word <= 'h0000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 84
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 332: ir 'h%h !== 'h0", ir); end	// Vector No: 83
assert (op === 'h00) else begin fail = 1; $display("Error 333: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 334: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 335: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000000000200000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000200000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 85
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 336: ir 'h%h !== 'h0", ir); end	// Vector No: 84
assert (op === 'h00) else begin fail = 1; $display("Error 337: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 338: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 339: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000200000:0:1:0:02:0:00000:
//------------------------

#2;
word <= 'h0000000000200000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 86
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 340: ir 'h%h !== 'h0", ir); end	// Vector No: 85
assert (op === 'h02) else begin fail = 1; $display("Error 341: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 342: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 343: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000200000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000200000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 87
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 344: ir 'h%h !== 'h0", ir); end	// Vector No: 86
assert (op === 'h00) else begin fail = 1; $display("Error 345: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 346: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 347: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000200000:1:1:0:00:0:00200:
//------------------------

#2;
word <= 'h0000000000200000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 88
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 348: ir 'h%h !== 'h0", ir); end	// Vector No: 87
assert (op === 'h00) else begin fail = 1; $display("Error 349: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 350: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 351: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000000000400000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000400000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 89
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 352: ir 'h%h !== 'h0", ir); end	// Vector No: 88
assert (op === 'h00) else begin fail = 1; $display("Error 353: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 354: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 355: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000400000:0:1:0:04:0:00000:
//------------------------

#2;
word <= 'h0000000000400000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 90
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 356: ir 'h%h !== 'h0", ir); end	// Vector No: 89
assert (op === 'h04) else begin fail = 1; $display("Error 357: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 358: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 359: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000400000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000400000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 91
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 360: ir 'h%h !== 'h0", ir); end	// Vector No: 90
assert (op === 'h00) else begin fail = 1; $display("Error 361: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 362: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 363: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000400000:1:1:0:00:0:00400:
//------------------------

#2;
word <= 'h0000000000400000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 92
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 364: ir 'h%h !== 'h0", ir); end	// Vector No: 91
assert (op === 'h00) else begin fail = 1; $display("Error 365: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 366: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 367: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000000000800000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000800000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 93
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 368: ir 'h%h !== 'h0", ir); end	// Vector No: 92
assert (op === 'h00) else begin fail = 1; $display("Error 369: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 370: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 371: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000800000:0:1:0:08:0:00000:
//------------------------

#2;
word <= 'h0000000000800000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 94
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 372: ir 'h%h !== 'h0", ir); end	// Vector No: 93
assert (op === 'h08) else begin fail = 1; $display("Error 373: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 374: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 375: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000800000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000000800000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 95
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 376: ir 'h%h !== 'h0", ir); end	// Vector No: 94
assert (op === 'h00) else begin fail = 1; $display("Error 377: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 378: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 379: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000000800000:1:1:0:00:0:00800:
//------------------------

#2;
word <= 'h0000000000800000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 96
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 380: ir 'h%h !== 'h0", ir); end	// Vector No: 95
assert (op === 'h00) else begin fail = 1; $display("Error 381: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 382: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 383: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000000001000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 97
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 384: ir 'h%h !== 'h0", ir); end	// Vector No: 96
assert (op === 'h00) else begin fail = 1; $display("Error 385: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 386: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 387: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000001000000:0:1:0:10:0:00000:
//------------------------

#2;
word <= 'h0000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 98
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 388: ir 'h%h !== 'h0", ir); end	// Vector No: 97
assert (op === 'h10) else begin fail = 1; $display("Error 389: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 390: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 391: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000001000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 99
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 392: ir 'h%h !== 'h0", ir); end	// Vector No: 98
assert (op === 'h00) else begin fail = 1; $display("Error 393: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 394: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 395: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000001000000:1:1:0:01:0:00000:
//------------------------

#2;
word <= 'h0000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 100
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 396: ir 'h%h !== 'h0", ir); end	// Vector No: 99
assert (op === 'h01) else begin fail = 1; $display("Error 397: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 398: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 399: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000002000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000002000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 101
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 400: ir 'h%h !== 'h0", ir); end	// Vector No: 100
assert (op === 'h00) else begin fail = 1; $display("Error 401: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 402: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 403: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000002000000:0:1:0:20:0:00000:
//------------------------

#2;
word <= 'h0000000002000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 102
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 404: ir 'h%h !== 'h0", ir); end	// Vector No: 101
assert (op === 'h20) else begin fail = 1; $display("Error 405: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 406: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 407: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000002000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000002000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 103
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 408: ir 'h%h !== 'h0", ir); end	// Vector No: 102
assert (op === 'h00) else begin fail = 1; $display("Error 409: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 410: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 411: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000002000000:1:1:0:02:0:00000:
//------------------------

#2;
word <= 'h0000000002000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 104
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 412: ir 'h%h !== 'h0", ir); end	// Vector No: 103
assert (op === 'h02) else begin fail = 1; $display("Error 413: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 414: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 415: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000004000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000004000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 105
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 416: ir 'h%h !== 'h0", ir); end	// Vector No: 104
assert (op === 'h00) else begin fail = 1; $display("Error 417: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 418: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 419: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000004000000:0:1:0:40:0:00000:
//------------------------

#2;
word <= 'h0000000004000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 106
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 420: ir 'h%h !== 'h0", ir); end	// Vector No: 105
assert (op === 'h40) else begin fail = 1; $display("Error 421: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 422: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 423: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000004000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000004000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 107
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 424: ir 'h%h !== 'h0", ir); end	// Vector No: 106
assert (op === 'h00) else begin fail = 1; $display("Error 425: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 426: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 427: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000004000000:1:1:0:04:0:00000:
//------------------------

#2;
word <= 'h0000000004000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 108
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 428: ir 'h%h !== 'h0", ir); end	// Vector No: 107
assert (op === 'h04) else begin fail = 1; $display("Error 429: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 430: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 431: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000008000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000008000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 109
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 432: ir 'h%h !== 'h0", ir); end	// Vector No: 108
assert (op === 'h00) else begin fail = 1; $display("Error 433: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 434: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 435: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000008000000:0:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000008000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 110
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 436: ir 'h%h !== 'h0", ir); end	// Vector No: 109
assert (op === 'h80) else begin fail = 1; $display("Error 437: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 438: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 439: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000008000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000008000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 111
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 440: ir 'h%h !== 'h0", ir); end	// Vector No: 110
assert (op === 'h00) else begin fail = 1; $display("Error 441: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 442: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 443: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000008000000:1:1:0:08:0:00000:
//------------------------

#2;
word <= 'h0000000008000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 112
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 444: ir 'h%h !== 'h0", ir); end	// Vector No: 111
assert (op === 'h08) else begin fail = 1; $display("Error 445: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 446: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 447: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000010000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 113
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 448: ir 'h%h !== 'h0", ir); end	// Vector No: 112
assert (op === 'h00) else begin fail = 1; $display("Error 449: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 450: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 451: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000010000000:0:1:1:00:0:00000:
//------------------------

#2;
word <= 'h0000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 114
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 452: ir 'h%h !== 'h1", ir); end	// Vector No: 113
assert (op === 'h00) else begin fail = 1; $display("Error 453: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 454: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 455: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000010000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 115
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 456: ir 'h%h !== 'h0", ir); end	// Vector No: 114
assert (op === 'h00) else begin fail = 1; $display("Error 457: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 458: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 459: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000010000000:1:1:0:10:0:00000:
//------------------------

#2;
word <= 'h0000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 116
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 460: ir 'h%h !== 'h0", ir); end	// Vector No: 115
assert (op === 'h10) else begin fail = 1; $display("Error 461: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 462: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 463: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000020000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000020000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 117
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 464: ir 'h%h !== 'h0", ir); end	// Vector No: 116
assert (op === 'h00) else begin fail = 1; $display("Error 465: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 466: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 467: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000020000000:0:1:2:00:0:00000:
//------------------------

#2;
word <= 'h0000000020000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 118
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 468: ir 'h%h !== 'h2", ir); end	// Vector No: 117
assert (op === 'h00) else begin fail = 1; $display("Error 469: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 470: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 471: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000020000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000020000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 119
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 472: ir 'h%h !== 'h0", ir); end	// Vector No: 118
assert (op === 'h00) else begin fail = 1; $display("Error 473: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 474: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 475: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000020000000:1:1:0:20:0:00000:
//------------------------

#2;
word <= 'h0000000020000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 120
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 476: ir 'h%h !== 'h0", ir); end	// Vector No: 119
assert (op === 'h20) else begin fail = 1; $display("Error 477: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 478: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 479: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000040000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000040000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 121
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 480: ir 'h%h !== 'h0", ir); end	// Vector No: 120
assert (op === 'h00) else begin fail = 1; $display("Error 481: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 482: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 483: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000040000000:0:1:4:00:0:00000:
//------------------------

#2;
word <= 'h0000000040000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 122
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 484: ir 'h%h !== 'h4", ir); end	// Vector No: 121
assert (op === 'h00) else begin fail = 1; $display("Error 485: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 486: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 487: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000040000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000040000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 123
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 488: ir 'h%h !== 'h0", ir); end	// Vector No: 122
assert (op === 'h00) else begin fail = 1; $display("Error 489: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 490: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 491: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000040000000:1:1:0:40:0:07000:
//------------------------

#2;
word <= 'h0000000040000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 124
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 492: ir 'h%h !== 'h0", ir); end	// Vector No: 123
assert (op === 'h40) else begin fail = 1; $display("Error 493: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 494: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 495: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0000000080000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 125
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 496: ir 'h%h !== 'h0", ir); end	// Vector No: 124
assert (op === 'h00) else begin fail = 1; $display("Error 497: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 498: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 499: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 126
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 500: ir 'h%h !== 'h8", ir); end	// Vector No: 125
assert (op === 'h00) else begin fail = 1; $display("Error 501: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 502: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 503: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 127
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 504: ir 'h%h !== 'h0", ir); end	// Vector No: 126
assert (op === 'h00) else begin fail = 1; $display("Error 505: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 506: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 507: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 128
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 508: ir 'h%h !== 'h0", ir); end	// Vector No: 127
assert (op === 'h80) else begin fail = 1; $display("Error 509: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 510: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 511: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000100000000:0:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 129
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 512: ir 'h%h !== 'h0", ir); end	// Vector No: 128
assert (op === 'h00) else begin fail = 1; $display("Error 513: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 514: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 515: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000100000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 130
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 516: ir 'h%h !== 'h0", ir); end	// Vector No: 129
assert (op === 'h00) else begin fail = 1; $display("Error 517: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 518: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 519: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000100000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 131
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 520: ir 'h%h !== 'h0", ir); end	// Vector No: 130
assert (op === 'h00) else begin fail = 1; $display("Error 521: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 522: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 523: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000100000000:1:1:1:00:0:00000:
//------------------------

#2;
word <= 'h0000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 132
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 524: ir 'h%h !== 'h1", ir); end	// Vector No: 131
assert (op === 'h00) else begin fail = 1; $display("Error 525: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 526: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 527: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000200000000:0:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000000200000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 133
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 528: ir 'h%h !== 'h0", ir); end	// Vector No: 132
assert (op === 'h00) else begin fail = 1; $display("Error 529: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 530: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 531: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000200000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000200000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 134
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 532: ir 'h%h !== 'h0", ir); end	// Vector No: 133
assert (op === 'h00) else begin fail = 1; $display("Error 533: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 534: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 535: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000200000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000200000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 135
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 536: ir 'h%h !== 'h0", ir); end	// Vector No: 134
assert (op === 'h00) else begin fail = 1; $display("Error 537: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 538: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 539: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000200000000:1:1:2:00:0:00000:
//------------------------

#2;
word <= 'h0000000200000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 136
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 540: ir 'h%h !== 'h2", ir); end	// Vector No: 135
assert (op === 'h00) else begin fail = 1; $display("Error 541: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 542: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 543: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000400000000:0:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000000400000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 137
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 544: ir 'h%h !== 'h0", ir); end	// Vector No: 136
assert (op === 'h00) else begin fail = 1; $display("Error 545: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 546: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 547: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000400000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000400000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 138
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 548: ir 'h%h !== 'h0", ir); end	// Vector No: 137
assert (op === 'h00) else begin fail = 1; $display("Error 549: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 550: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 551: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000400000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000400000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 139
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 552: ir 'h%h !== 'h0", ir); end	// Vector No: 138
assert (op === 'h00) else begin fail = 1; $display("Error 553: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 554: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 555: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000400000000:1:1:4:00:0:00000:
//------------------------

#2;
word <= 'h0000000400000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 140
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 556: ir 'h%h !== 'h4", ir); end	// Vector No: 139
assert (op === 'h00) else begin fail = 1; $display("Error 557: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 558: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 559: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000800000000:0:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000000800000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 141
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 560: ir 'h%h !== 'h0", ir); end	// Vector No: 140
assert (op === 'h00) else begin fail = 1; $display("Error 561: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 562: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 563: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000800000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000800000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 142
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 564: ir 'h%h !== 'h0", ir); end	// Vector No: 141
assert (op === 'h00) else begin fail = 1; $display("Error 565: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 566: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 567: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000800000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000800000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 143
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 568: ir 'h%h !== 'h0", ir); end	// Vector No: 142
assert (op === 'h00) else begin fail = 1; $display("Error 569: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 570: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 571: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000800000000:1:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000800000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 144
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 572: ir 'h%h !== 'h8", ir); end	// Vector No: 143
assert (op === 'h00) else begin fail = 1; $display("Error 573: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 574: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 575: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001000000000:0:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 145
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 576: ir 'h%h !== 'h0", ir); end	// Vector No: 144
assert (op === 'h00) else begin fail = 1; $display("Error 577: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 578: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 579: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000001000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 146
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 580: ir 'h%h !== 'h0", ir); end	// Vector No: 145
assert (op === 'h00) else begin fail = 1; $display("Error 581: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 582: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 583: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001000000000:1:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 147
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 584: ir 'h%h !== 'h0", ir); end	// Vector No: 146
assert (op === 'h00) else begin fail = 1; $display("Error 585: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 586: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 587: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000001000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 148
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 588: ir 'h%h !== 'h0", ir); end	// Vector No: 147
assert (op === 'h00) else begin fail = 1; $display("Error 589: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 590: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 591: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002000000000:0:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000002000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 149
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 592: ir 'h%h !== 'h0", ir); end	// Vector No: 148
assert (op === 'h00) else begin fail = 1; $display("Error 593: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 594: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 595: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000002000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000002000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 150
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 596: ir 'h%h !== 'h0", ir); end	// Vector No: 149
assert (op === 'h00) else begin fail = 1; $display("Error 597: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 598: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 599: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002000000000:1:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000002000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 151
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 600: ir 'h%h !== 'h0", ir); end	// Vector No: 150
assert (op === 'h00) else begin fail = 1; $display("Error 601: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 602: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 603: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000002000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000002000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 152
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 604: ir 'h%h !== 'h0", ir); end	// Vector No: 151
assert (op === 'h00) else begin fail = 1; $display("Error 605: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 606: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 607: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004000000000:0:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000004000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 153
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 608: ir 'h%h !== 'h0", ir); end	// Vector No: 152
assert (op === 'h00) else begin fail = 1; $display("Error 609: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 610: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 611: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000004000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000004000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 154
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 612: ir 'h%h !== 'h0", ir); end	// Vector No: 153
assert (op === 'h00) else begin fail = 1; $display("Error 613: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 614: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 615: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004000000000:1:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000004000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 155
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 616: ir 'h%h !== 'h0", ir); end	// Vector No: 154
assert (op === 'h00) else begin fail = 1; $display("Error 617: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 618: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 619: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000004000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000004000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 156
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 620: ir 'h%h !== 'h0", ir); end	// Vector No: 155
assert (op === 'h00) else begin fail = 1; $display("Error 621: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 622: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 623: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008000000000:0:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000008000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 157
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 624: ir 'h%h !== 'h0", ir); end	// Vector No: 156
assert (op === 'h00) else begin fail = 1; $display("Error 625: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 626: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 627: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000008000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000008000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 158
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 628: ir 'h%h !== 'h0", ir); end	// Vector No: 157
assert (op === 'h00) else begin fail = 1; $display("Error 629: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 630: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 631: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008000000000:1:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000008000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 159
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 632: ir 'h%h !== 'h0", ir); end	// Vector No: 158
assert (op === 'h00) else begin fail = 1; $display("Error 633: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 634: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 635: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000008000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000008000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 160
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 636: ir 'h%h !== 'h0", ir); end	// Vector No: 159
assert (op === 'h00) else begin fail = 1; $display("Error 637: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 638: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 639: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010000000000:0:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 161
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 640: ir 'h%h !== 'h0", ir); end	// Vector No: 160
assert (op === 'h00) else begin fail = 1; $display("Error 641: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 642: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 643: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000010000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 162
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 644: ir 'h%h !== 'h0", ir); end	// Vector No: 161
assert (op === 'h00) else begin fail = 1; $display("Error 645: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 646: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 647: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010000000000:1:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 163
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 648: ir 'h%h !== 'h0", ir); end	// Vector No: 162
assert (op === 'h00) else begin fail = 1; $display("Error 649: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 650: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 651: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000010000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 164
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 652: ir 'h%h !== 'h0", ir); end	// Vector No: 163
assert (op === 'h00) else begin fail = 1; $display("Error 653: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 654: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 655: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020000000000:0:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000020000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 165
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 656: ir 'h%h !== 'h0", ir); end	// Vector No: 164
assert (op === 'h00) else begin fail = 1; $display("Error 657: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 658: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 659: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000020000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000020000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 166
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 660: ir 'h%h !== 'h0", ir); end	// Vector No: 165
assert (op === 'h00) else begin fail = 1; $display("Error 661: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 662: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 663: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020000000000:1:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000020000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 167
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 664: ir 'h%h !== 'h0", ir); end	// Vector No: 166
assert (op === 'h00) else begin fail = 1; $display("Error 665: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 666: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 667: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000020000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000020000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 168
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 668: ir 'h%h !== 'h0", ir); end	// Vector No: 167
assert (op === 'h00) else begin fail = 1; $display("Error 669: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 670: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 671: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040000000000:0:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000040000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 169
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 672: ir 'h%h !== 'h0", ir); end	// Vector No: 168
assert (op === 'h00) else begin fail = 1; $display("Error 673: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 674: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 675: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000040000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000040000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 170
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 676: ir 'h%h !== 'h0", ir); end	// Vector No: 169
assert (op === 'h00) else begin fail = 1; $display("Error 677: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 678: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 679: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040000000000:1:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000040000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 171
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 680: ir 'h%h !== 'h0", ir); end	// Vector No: 170
assert (op === 'h00) else begin fail = 1; $display("Error 681: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 682: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 683: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000040000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000040000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 172
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 684: ir 'h%h !== 'h0", ir); end	// Vector No: 171
assert (op === 'h00) else begin fail = 1; $display("Error 685: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 686: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 687: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080000000000:0:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000080000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 173
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 688: ir 'h%h !== 'h0", ir); end	// Vector No: 172
assert (op === 'h00) else begin fail = 1; $display("Error 689: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 690: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 691: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000080000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000080000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 174
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 692: ir 'h%h !== 'h0", ir); end	// Vector No: 173
assert (op === 'h00) else begin fail = 1; $display("Error 693: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 694: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 695: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080000000000:1:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000080000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 175
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 696: ir 'h%h !== 'h0", ir); end	// Vector No: 174
assert (op === 'h00) else begin fail = 1; $display("Error 697: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 698: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 699: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000080000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000080000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 176
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 700: ir 'h%h !== 'h0", ir); end	// Vector No: 175
assert (op === 'h00) else begin fail = 1; $display("Error 701: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 702: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 703: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100000000000:0:0:0:00:0:01000:
//------------------------

#2;
word <= 'h0000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 177
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 704: ir 'h%h !== 'h0", ir); end	// Vector No: 176
assert (op === 'h00) else begin fail = 1; $display("Error 705: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 706: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 707: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000100000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 178
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 708: ir 'h%h !== 'h0", ir); end	// Vector No: 177
assert (op === 'h00) else begin fail = 1; $display("Error 709: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 710: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 711: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100000000000:1:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 179
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 712: ir 'h%h !== 'h0", ir); end	// Vector No: 178
assert (op === 'h00) else begin fail = 1; $display("Error 713: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 714: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 715: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000100000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 180
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 716: ir 'h%h !== 'h0", ir); end	// Vector No: 179
assert (op === 'h00) else begin fail = 1; $display("Error 717: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 718: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 719: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200000000000:0:0:0:00:0:02000:
//------------------------

#2;
word <= 'h0000200000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 181
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 720: ir 'h%h !== 'h0", ir); end	// Vector No: 180
assert (op === 'h00) else begin fail = 1; $display("Error 721: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 722: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 723: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000200000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000200000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 182
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 724: ir 'h%h !== 'h0", ir); end	// Vector No: 181
assert (op === 'h00) else begin fail = 1; $display("Error 725: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 726: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 727: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200000000000:1:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000200000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 183
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 728: ir 'h%h !== 'h0", ir); end	// Vector No: 182
assert (op === 'h00) else begin fail = 1; $display("Error 729: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 730: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 731: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000200000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000200000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 184
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 732: ir 'h%h !== 'h0", ir); end	// Vector No: 183
assert (op === 'h00) else begin fail = 1; $display("Error 733: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 734: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 735: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400000000000:0:0:0:00:0:04000:
//------------------------

#2;
word <= 'h0000400000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 185
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 736: ir 'h%h !== 'h0", ir); end	// Vector No: 184
assert (op === 'h00) else begin fail = 1; $display("Error 737: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 738: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 739: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000400000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000400000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 186
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 740: ir 'h%h !== 'h0", ir); end	// Vector No: 185
assert (op === 'h00) else begin fail = 1; $display("Error 741: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 742: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 743: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400000000000:1:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000400000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 187
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 744: ir 'h%h !== 'h0", ir); end	// Vector No: 186
assert (op === 'h00) else begin fail = 1; $display("Error 745: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 746: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 747: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000400000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000400000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 188
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 748: ir 'h%h !== 'h0", ir); end	// Vector No: 187
assert (op === 'h00) else begin fail = 1; $display("Error 749: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 750: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 751: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800000000000:0:0:0:00:0:08000:
//------------------------

#2;
word <= 'h0000800000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 189
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 752: ir 'h%h !== 'h0", ir); end	// Vector No: 188
assert (op === 'h00) else begin fail = 1; $display("Error 753: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 754: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 755: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000800000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000800000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 190
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 756: ir 'h%h !== 'h0", ir); end	// Vector No: 189
assert (op === 'h00) else begin fail = 1; $display("Error 757: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 758: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 759: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800000000000:1:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000800000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 191
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 760: ir 'h%h !== 'h0", ir); end	// Vector No: 190
assert (op === 'h00) else begin fail = 1; $display("Error 761: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 762: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 763: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000800000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0000800000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 192
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 764: ir 'h%h !== 'h0", ir); end	// Vector No: 191
assert (op === 'h00) else begin fail = 1; $display("Error 765: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 766: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 767: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000000000000:0:0:0:00:0:10000:
//------------------------

#2;
word <= 'h0001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 193
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 768: ir 'h%h !== 'h0", ir); end	// Vector No: 192
assert (op === 'h00) else begin fail = 1; $display("Error 769: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 770: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 771: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0001000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 194
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 772: ir 'h%h !== 'h0", ir); end	// Vector No: 193
assert (op === 'h00) else begin fail = 1; $display("Error 773: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 774: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 775: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000000000000:1:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 195
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 776: ir 'h%h !== 'h0", ir); end	// Vector No: 194
assert (op === 'h01) else begin fail = 1; $display("Error 777: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 778: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 779: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 196
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 780: ir 'h%h !== 'h0", ir); end	// Vector No: 195
assert (op === 'h00) else begin fail = 1; $display("Error 781: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 782: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 783: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000000000000:0:0:0:00:0:20000:
//------------------------

#2;
word <= 'h0002000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 197
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 784: ir 'h%h !== 'h0", ir); end	// Vector No: 196
assert (op === 'h00) else begin fail = 1; $display("Error 785: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 786: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 787: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0002000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0002000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 198
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 788: ir 'h%h !== 'h0", ir); end	// Vector No: 197
assert (op === 'h00) else begin fail = 1; $display("Error 789: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 790: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 791: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000000000000:1:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0002000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 199
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 792: ir 'h%h !== 'h0", ir); end	// Vector No: 198
assert (op === 'h02) else begin fail = 1; $display("Error 793: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 794: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 795: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0002000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 200
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 796: ir 'h%h !== 'h0", ir); end	// Vector No: 199
assert (op === 'h00) else begin fail = 1; $display("Error 797: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 798: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 799: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000000000000:0:0:0:00:0:40000:
//------------------------

#2;
word <= 'h0004000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 201
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 800: ir 'h%h !== 'h0", ir); end	// Vector No: 200
assert (op === 'h00) else begin fail = 1; $display("Error 801: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 802: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 803: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0004000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0004000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 202
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 804: ir 'h%h !== 'h0", ir); end	// Vector No: 201
assert (op === 'h00) else begin fail = 1; $display("Error 805: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 806: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 807: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000000000000:1:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0004000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 203
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 808: ir 'h%h !== 'h0", ir); end	// Vector No: 202
assert (op === 'h04) else begin fail = 1; $display("Error 809: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 810: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 811: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0004000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 204
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 812: ir 'h%h !== 'h0", ir); end	// Vector No: 203
assert (op === 'h00) else begin fail = 1; $display("Error 813: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 814: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 815: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000000000000:0:0:0:00:0:80000:
//------------------------

#2;
word <= 'h0008000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 205
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 816: ir 'h%h !== 'h0", ir); end	// Vector No: 204
assert (op === 'h00) else begin fail = 1; $display("Error 817: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 818: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 819: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0008000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0008000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 206
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 820: ir 'h%h !== 'h0", ir); end	// Vector No: 205
assert (op === 'h00) else begin fail = 1; $display("Error 821: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 822: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 823: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000000000000:1:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0008000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 207
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 824: ir 'h%h !== 'h0", ir); end	// Vector No: 206
assert (op === 'h08) else begin fail = 1; $display("Error 825: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 826: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 827: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0008000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 208
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 828: ir 'h%h !== 'h0", ir); end	// Vector No: 207
assert (op === 'h00) else begin fail = 1; $display("Error 829: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 830: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 831: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000000000000:0:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 209
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 832: ir 'h%h !== 'h0", ir); end	// Vector No: 208
assert (op === 'h01) else begin fail = 1; $display("Error 833: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 834: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 835: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 210
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 836: ir 'h%h !== 'h0", ir); end	// Vector No: 209
assert (op === 'h00) else begin fail = 1; $display("Error 837: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 838: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 839: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000000000000:1:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 211
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 840: ir 'h%h !== 'h0", ir); end	// Vector No: 210
assert (op === 'h10) else begin fail = 1; $display("Error 841: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 842: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 843: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 212
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 844: ir 'h%h !== 'h0", ir); end	// Vector No: 211
assert (op === 'h00) else begin fail = 1; $display("Error 845: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 846: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 847: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000000000000:0:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0020000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 213
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 848: ir 'h%h !== 'h0", ir); end	// Vector No: 212
assert (op === 'h02) else begin fail = 1; $display("Error 849: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 850: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 851: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0020000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 214
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 852: ir 'h%h !== 'h0", ir); end	// Vector No: 213
assert (op === 'h00) else begin fail = 1; $display("Error 853: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 854: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 855: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000000000000:1:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0020000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 215
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 856: ir 'h%h !== 'h0", ir); end	// Vector No: 214
assert (op === 'h20) else begin fail = 1; $display("Error 857: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 858: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 859: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0020000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 216
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 860: ir 'h%h !== 'h0", ir); end	// Vector No: 215
assert (op === 'h00) else begin fail = 1; $display("Error 861: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 862: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 863: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000000000000:0:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0040000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 217
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 864: ir 'h%h !== 'h0", ir); end	// Vector No: 216
assert (op === 'h04) else begin fail = 1; $display("Error 865: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 866: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 867: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0040000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 218
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 868: ir 'h%h !== 'h0", ir); end	// Vector No: 217
assert (op === 'h00) else begin fail = 1; $display("Error 869: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 870: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 871: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000000000000:1:0:0:40:0:07000:
//------------------------

#2;
word <= 'h0040000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 219
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 872: ir 'h%h !== 'h0", ir); end	// Vector No: 218
assert (op === 'h40) else begin fail = 1; $display("Error 873: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 874: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 875: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0040000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0040000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 220
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 876: ir 'h%h !== 'h0", ir); end	// Vector No: 219
assert (op === 'h00) else begin fail = 1; $display("Error 877: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 878: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 879: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 221
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 880: ir 'h%h !== 'h0", ir); end	// Vector No: 220
assert (op === 'h08) else begin fail = 1; $display("Error 881: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 882: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 883: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 222
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 884: ir 'h%h !== 'h0", ir); end	// Vector No: 221
assert (op === 'h00) else begin fail = 1; $display("Error 885: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 886: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 887: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 223
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 888: ir 'h%h !== 'h0", ir); end	// Vector No: 222
assert (op === 'h80) else begin fail = 1; $display("Error 889: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 890: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 891: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 224
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 892: ir 'h%h !== 'h0", ir); end	// Vector No: 223
assert (op === 'h00) else begin fail = 1; $display("Error 893: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 894: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 895: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000000000000:0:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 225
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 896: ir 'h%h !== 'h0", ir); end	// Vector No: 224
assert (op === 'h10) else begin fail = 1; $display("Error 897: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 898: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 899: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 226
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 900: ir 'h%h !== 'h0", ir); end	// Vector No: 225
assert (op === 'h00) else begin fail = 1; $display("Error 901: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 902: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 903: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000000000000:1:0:1:00:0:00000:
//------------------------

#2;
word <= 'h0100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 227
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 904: ir 'h%h !== 'h1", ir); end	// Vector No: 226
assert (op === 'h00) else begin fail = 1; $display("Error 905: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 906: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 907: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 228
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 908: ir 'h%h !== 'h0", ir); end	// Vector No: 227
assert (op === 'h00) else begin fail = 1; $display("Error 909: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 910: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 911: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000000000000:0:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0200000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 229
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 912: ir 'h%h !== 'h0", ir); end	// Vector No: 228
assert (op === 'h20) else begin fail = 1; $display("Error 913: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 914: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 915: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0200000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 230
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 916: ir 'h%h !== 'h0", ir); end	// Vector No: 229
assert (op === 'h00) else begin fail = 1; $display("Error 917: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 918: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 919: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000000000000:1:0:2:00:0:00000:
//------------------------

#2;
word <= 'h0200000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 231
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 920: ir 'h%h !== 'h2", ir); end	// Vector No: 230
assert (op === 'h00) else begin fail = 1; $display("Error 921: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 922: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 923: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0200000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 232
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 924: ir 'h%h !== 'h0", ir); end	// Vector No: 231
assert (op === 'h00) else begin fail = 1; $display("Error 925: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 926: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 927: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000000000000:0:0:0:40:0:00000:
//------------------------

#2;
word <= 'h0400000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 233
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 928: ir 'h%h !== 'h0", ir); end	// Vector No: 232
assert (op === 'h40) else begin fail = 1; $display("Error 929: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 930: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 931: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0400000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 234
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 932: ir 'h%h !== 'h0", ir); end	// Vector No: 233
assert (op === 'h00) else begin fail = 1; $display("Error 933: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 934: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 935: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000000000000:1:0:4:00:0:00000:
//------------------------

#2;
word <= 'h0400000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 235
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 936: ir 'h%h !== 'h4", ir); end	// Vector No: 234
assert (op === 'h00) else begin fail = 1; $display("Error 937: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 938: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 939: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0400000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 236
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 940: ir 'h%h !== 'h0", ir); end	// Vector No: 235
assert (op === 'h00) else begin fail = 1; $display("Error 941: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 942: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 943: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000000000000:0:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0800000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 237
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 944: ir 'h%h !== 'h0", ir); end	// Vector No: 236
assert (op === 'h80) else begin fail = 1; $display("Error 945: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 946: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 947: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0800000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 238
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 948: ir 'h%h !== 'h0", ir); end	// Vector No: 237
assert (op === 'h00) else begin fail = 1; $display("Error 949: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 950: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 951: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000000000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0800000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 239
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 952: ir 'h%h !== 'h0", ir); end	// Vector No: 238
assert (op === 'h00) else begin fail = 1; $display("Error 953: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 954: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 955: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0800000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 240
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 956: ir 'h%h !== 'h0", ir); end	// Vector No: 239
assert (op === 'h00) else begin fail = 1; $display("Error 957: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 958: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 959: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000000000000:0:0:1:00:0:00000:
//------------------------

#2;
word <= 'h1000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 241
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 960: ir 'h%h !== 'h1", ir); end	// Vector No: 240
assert (op === 'h00) else begin fail = 1; $display("Error 961: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 962: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 963: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h1000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 242
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 964: ir 'h%h !== 'h0", ir); end	// Vector No: 241
assert (op === 'h00) else begin fail = 1; $display("Error 965: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 966: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 967: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000000000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h1000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 243
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 968: ir 'h%h !== 'h0", ir); end	// Vector No: 242
assert (op === 'h00) else begin fail = 1; $display("Error 969: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 970: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 971: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h1000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 244
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 972: ir 'h%h !== 'h0", ir); end	// Vector No: 243
assert (op === 'h00) else begin fail = 1; $display("Error 973: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 974: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 975: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000000000000:0:0:2:00:0:00000:
//------------------------

#2;
word <= 'h2000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 245
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 976: ir 'h%h !== 'h2", ir); end	// Vector No: 244
assert (op === 'h00) else begin fail = 1; $display("Error 977: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 978: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 979: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h2000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 246
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 980: ir 'h%h !== 'h0", ir); end	// Vector No: 245
assert (op === 'h00) else begin fail = 1; $display("Error 981: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 982: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 983: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000000000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h2000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 247
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 984: ir 'h%h !== 'h0", ir); end	// Vector No: 246
assert (op === 'h00) else begin fail = 1; $display("Error 985: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 986: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 987: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h2000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 248
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 988: ir 'h%h !== 'h0", ir); end	// Vector No: 247
assert (op === 'h00) else begin fail = 1; $display("Error 989: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 990: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 991: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000000000000:0:0:4:00:0:00000:
//------------------------

#2;
word <= 'h4000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 249
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 992: ir 'h%h !== 'h4", ir); end	// Vector No: 248
assert (op === 'h00) else begin fail = 1; $display("Error 993: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 994: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 995: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h4000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 250
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 996: ir 'h%h !== 'h0", ir); end	// Vector No: 249
assert (op === 'h00) else begin fail = 1; $display("Error 997: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 998: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 999: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000000000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h4000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 251
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 1000: ir 'h%h !== 'h0", ir); end	// Vector No: 250
assert (op === 'h00) else begin fail = 1; $display("Error 1001: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1002: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1003: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h4000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 252
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 1004: ir 'h%h !== 'h0", ir); end	// Vector No: 251
assert (op === 'h00) else begin fail = 1; $display("Error 1005: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1006: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1007: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000000000000:0:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 253
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 1008: ir 'h%h !== 'h8", ir); end	// Vector No: 252
assert (op === 'h00) else begin fail = 1; $display("Error 1009: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1010: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1011: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h8000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 254
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 1012: ir 'h%h !== 'h0", ir); end	// Vector No: 253
assert (op === 'h00) else begin fail = 1; $display("Error 1013: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1014: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1015: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000000000000:1:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 255
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 1016: ir 'h%h !== 'h8", ir); end	// Vector No: 254
assert (op === 'h00) else begin fail = 1; $display("Error 1017: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1018: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1019: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h8000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 256
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 1020: ir 'h%h !== 'h0", ir); end	// Vector No: 255
assert (op === 'h00) else begin fail = 1; $display("Error 1021: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1022: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 1023: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// fffffffffffffffe:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffffe;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 257
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1024: ir 'h%h !== 'hf", ir); end	// Vector No: 256
assert (op === 'hff) else begin fail = 1; $display("Error 1025: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1026: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1027: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffffe:0:1:f:ff:0:ffffe:
//------------------------

#2;
word <= 'hfffffffffffffffe;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 258
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1028: ir 'h%h !== 'hf", ir); end	// Vector No: 257
assert (op === 'hff) else begin fail = 1; $display("Error 1029: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1030: extop 'h%h !== 0", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 1031: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// fffffffffffffffe:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffe;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 259
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1032: ir 'h%h !== 'hf", ir); end	// Vector No: 258
assert (op === 'hf8) else begin fail = 1; $display("Error 1033: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1034: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1035: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffffe:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffe;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 260
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1036: ir 'h%h !== 'hf", ir); end	// Vector No: 259
assert (op === 'hf8) else begin fail = 1; $display("Error 1037: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1038: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1039: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffffd:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffffd;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 261
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1040: ir 'h%h !== 'hf", ir); end	// Vector No: 260
assert (op === 'hff) else begin fail = 1; $display("Error 1041: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1042: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1043: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffffd:0:1:f:ff:0:ffffd:
//------------------------

#2;
word <= 'hfffffffffffffffd;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 262
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1044: ir 'h%h !== 'hf", ir); end	// Vector No: 261
assert (op === 'hff) else begin fail = 1; $display("Error 1045: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1046: extop 'h%h !== 0", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 1047: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// fffffffffffffffd:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffd;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 263
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1048: ir 'h%h !== 'hf", ir); end	// Vector No: 262
assert (op === 'hf8) else begin fail = 1; $display("Error 1049: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1050: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1051: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffffd:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffd;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 264
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1052: ir 'h%h !== 'hf", ir); end	// Vector No: 263
assert (op === 'hf8) else begin fail = 1; $display("Error 1053: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1054: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1055: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffffb:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffffb;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 265
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1056: ir 'h%h !== 'hf", ir); end	// Vector No: 264
assert (op === 'hff) else begin fail = 1; $display("Error 1057: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1058: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1059: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffffb:0:1:f:ff:0:ffffb:
//------------------------

#2;
word <= 'hfffffffffffffffb;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 266
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1060: ir 'h%h !== 'hf", ir); end	// Vector No: 265
assert (op === 'hff) else begin fail = 1; $display("Error 1061: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1062: extop 'h%h !== 0", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 1063: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// fffffffffffffffb:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffb;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 267
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1064: ir 'h%h !== 'hf", ir); end	// Vector No: 266
assert (op === 'hf8) else begin fail = 1; $display("Error 1065: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1066: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1067: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffffb:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffffb;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 268
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1068: ir 'h%h !== 'hf", ir); end	// Vector No: 267
assert (op === 'hf8) else begin fail = 1; $display("Error 1069: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1070: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1071: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffff7:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffff7;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 269
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1072: ir 'h%h !== 'hf", ir); end	// Vector No: 268
assert (op === 'hff) else begin fail = 1; $display("Error 1073: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1074: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1075: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffff7:0:1:f:ff:0:ffff7:
//------------------------

#2;
word <= 'hfffffffffffffff7;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 270
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1076: ir 'h%h !== 'hf", ir); end	// Vector No: 269
assert (op === 'hff) else begin fail = 1; $display("Error 1077: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1078: extop 'h%h !== 0", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 1079: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// fffffffffffffff7:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffff7;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 271
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1080: ir 'h%h !== 'hf", ir); end	// Vector No: 270
assert (op === 'hf8) else begin fail = 1; $display("Error 1081: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1082: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1083: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffff7:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffff7;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 272
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1084: ir 'h%h !== 'hf", ir); end	// Vector No: 271
assert (op === 'hf8) else begin fail = 1; $display("Error 1085: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1086: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1087: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffef:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffffef;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 273
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1088: ir 'h%h !== 'hf", ir); end	// Vector No: 272
assert (op === 'hff) else begin fail = 1; $display("Error 1089: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1090: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1091: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffffef:0:1:f:ff:0:fffef:
//------------------------

#2;
word <= 'hffffffffffffffef;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 274
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1092: ir 'h%h !== 'hf", ir); end	// Vector No: 273
assert (op === 'hff) else begin fail = 1; $display("Error 1093: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1094: extop 'h%h !== 0", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 1095: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// ffffffffffffffef:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffef;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 275
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1096: ir 'h%h !== 'hf", ir); end	// Vector No: 274
assert (op === 'hf8) else begin fail = 1; $display("Error 1097: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1098: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1099: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffef:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffef;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 276
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1100: ir 'h%h !== 'hf", ir); end	// Vector No: 275
assert (op === 'hf8) else begin fail = 1; $display("Error 1101: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1102: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1103: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffdf:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffffdf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 277
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1104: ir 'h%h !== 'hf", ir); end	// Vector No: 276
assert (op === 'hff) else begin fail = 1; $display("Error 1105: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1106: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1107: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffffdf:0:1:f:ff:0:fffdf:
//------------------------

#2;
word <= 'hffffffffffffffdf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 278
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1108: ir 'h%h !== 'hf", ir); end	// Vector No: 277
assert (op === 'hff) else begin fail = 1; $display("Error 1109: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1110: extop 'h%h !== 0", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 1111: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// ffffffffffffffdf:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffdf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 279
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1112: ir 'h%h !== 'hf", ir); end	// Vector No: 278
assert (op === 'hf8) else begin fail = 1; $display("Error 1113: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1114: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1115: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffdf:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffdf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 280
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1116: ir 'h%h !== 'hf", ir); end	// Vector No: 279
assert (op === 'hf8) else begin fail = 1; $display("Error 1117: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1118: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1119: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffbf:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffffbf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 281
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1120: ir 'h%h !== 'hf", ir); end	// Vector No: 280
assert (op === 'hff) else begin fail = 1; $display("Error 1121: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1122: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1123: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffffbf:0:1:f:ff:0:fffbf:
//------------------------

#2;
word <= 'hffffffffffffffbf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 282
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1124: ir 'h%h !== 'hf", ir); end	// Vector No: 281
assert (op === 'hff) else begin fail = 1; $display("Error 1125: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1126: extop 'h%h !== 0", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 1127: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// ffffffffffffffbf:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffbf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 283
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1128: ir 'h%h !== 'hf", ir); end	// Vector No: 282
assert (op === 'hf8) else begin fail = 1; $display("Error 1129: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1130: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1131: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffffbf:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffffbf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 284
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1132: ir 'h%h !== 'hf", ir); end	// Vector No: 283
assert (op === 'hf8) else begin fail = 1; $display("Error 1133: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1134: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1135: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffff7f:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffff7f;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 285
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1136: ir 'h%h !== 'hf", ir); end	// Vector No: 284
assert (op === 'hff) else begin fail = 1; $display("Error 1137: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1138: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1139: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffff7f:0:1:f:ff:0:fff7f:
//------------------------

#2;
word <= 'hffffffffffffff7f;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 286
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1140: ir 'h%h !== 'hf", ir); end	// Vector No: 285
assert (op === 'hff) else begin fail = 1; $display("Error 1141: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1142: extop 'h%h !== 0", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 1143: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// ffffffffffffff7f:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffff7f;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 287
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1144: ir 'h%h !== 'hf", ir); end	// Vector No: 286
assert (op === 'hf8) else begin fail = 1; $display("Error 1145: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1146: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1147: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffff7f:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffff7f;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 288
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1148: ir 'h%h !== 'hf", ir); end	// Vector No: 287
assert (op === 'hf8) else begin fail = 1; $display("Error 1149: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1150: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1151: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffeff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffeff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 289
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1152: ir 'h%h !== 'hf", ir); end	// Vector No: 288
assert (op === 'hff) else begin fail = 1; $display("Error 1153: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1154: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1155: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffeff:0:1:f:ff:0:ffeff:
//------------------------

#2;
word <= 'hfffffffffffffeff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 290
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1156: ir 'h%h !== 'hf", ir); end	// Vector No: 289
assert (op === 'hff) else begin fail = 1; $display("Error 1157: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1158: extop 'h%h !== 0", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 1159: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// fffffffffffffeff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffeff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 291
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1160: ir 'h%h !== 'hf", ir); end	// Vector No: 290
assert (op === 'hf8) else begin fail = 1; $display("Error 1161: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1162: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1163: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffeff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffeff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 292
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1164: ir 'h%h !== 'hf", ir); end	// Vector No: 291
assert (op === 'hf8) else begin fail = 1; $display("Error 1165: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1166: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1167: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffdff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffdff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 293
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1168: ir 'h%h !== 'hf", ir); end	// Vector No: 292
assert (op === 'hff) else begin fail = 1; $display("Error 1169: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1170: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1171: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffdff:0:1:f:ff:0:ffdff:
//------------------------

#2;
word <= 'hfffffffffffffdff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 294
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1172: ir 'h%h !== 'hf", ir); end	// Vector No: 293
assert (op === 'hff) else begin fail = 1; $display("Error 1173: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1174: extop 'h%h !== 0", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 1175: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// fffffffffffffdff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffdff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 295
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1176: ir 'h%h !== 'hf", ir); end	// Vector No: 294
assert (op === 'hf8) else begin fail = 1; $display("Error 1177: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1178: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1179: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffdff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffdff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 296
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1180: ir 'h%h !== 'hf", ir); end	// Vector No: 295
assert (op === 'hf8) else begin fail = 1; $display("Error 1181: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1182: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1183: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffbff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffffbff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 297
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1184: ir 'h%h !== 'hf", ir); end	// Vector No: 296
assert (op === 'hff) else begin fail = 1; $display("Error 1185: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1186: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1187: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffffbff:0:1:f:ff:0:ffbff:
//------------------------

#2;
word <= 'hfffffffffffffbff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 298
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1188: ir 'h%h !== 'hf", ir); end	// Vector No: 297
assert (op === 'hff) else begin fail = 1; $display("Error 1189: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1190: extop 'h%h !== 0", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 1191: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// fffffffffffffbff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffbff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 299
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1192: ir 'h%h !== 'hf", ir); end	// Vector No: 298
assert (op === 'hf8) else begin fail = 1; $display("Error 1193: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1194: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1195: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffffbff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffffbff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 300
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1196: ir 'h%h !== 'hf", ir); end	// Vector No: 299
assert (op === 'hf8) else begin fail = 1; $display("Error 1197: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1198: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1199: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffff7ff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffff7ff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 301
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1200: ir 'h%h !== 'hf", ir); end	// Vector No: 300
assert (op === 'hff) else begin fail = 1; $display("Error 1201: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1202: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1203: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffff7ff:0:1:f:ff:0:ff7ff:
//------------------------

#2;
word <= 'hfffffffffffff7ff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 302
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1204: ir 'h%h !== 'hf", ir); end	// Vector No: 301
assert (op === 'hff) else begin fail = 1; $display("Error 1205: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1206: extop 'h%h !== 0", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 1207: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// fffffffffffff7ff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffff7ff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 303
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1208: ir 'h%h !== 'hf", ir); end	// Vector No: 302
assert (op === 'hf8) else begin fail = 1; $display("Error 1209: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1210: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1211: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffff7ff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffff7ff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 304
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1212: ir 'h%h !== 'hf", ir); end	// Vector No: 303
assert (op === 'hf8) else begin fail = 1; $display("Error 1213: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1214: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1215: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffefff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffefff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 305
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1216: ir 'h%h !== 'hf", ir); end	// Vector No: 304
assert (op === 'hff) else begin fail = 1; $display("Error 1217: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1218: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1219: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffefff:0:1:f:ff:0:fefff:
//------------------------

#2;
word <= 'hffffffffffffefff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 306
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1220: ir 'h%h !== 'hf", ir); end	// Vector No: 305
assert (op === 'hff) else begin fail = 1; $display("Error 1221: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1222: extop 'h%h !== 0", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 1223: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// ffffffffffffefff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffefff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 307
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1224: ir 'h%h !== 'hf", ir); end	// Vector No: 306
assert (op === 'hf8) else begin fail = 1; $display("Error 1225: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1226: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1227: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffefff:1:1:f:f8:0:07ffe:
//------------------------

#2;
word <= 'hffffffffffffefff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 308
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1228: ir 'h%h !== 'hf", ir); end	// Vector No: 307
assert (op === 'hf8) else begin fail = 1; $display("Error 1229: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1230: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffe) else begin fail = 1; $display("Error 1231: addr 'h%h !== 'h07ffe", addr); end
#2;
clk <= 0;

// ffffffffffffdfff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffdfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 309
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1232: ir 'h%h !== 'hf", ir); end	// Vector No: 308
assert (op === 'hff) else begin fail = 1; $display("Error 1233: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1234: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1235: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffdfff:0:1:f:ff:0:fdfff:
//------------------------

#2;
word <= 'hffffffffffffdfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 310
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1236: ir 'h%h !== 'hf", ir); end	// Vector No: 309
assert (op === 'hff) else begin fail = 1; $display("Error 1237: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1238: extop 'h%h !== 0", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 1239: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// ffffffffffffdfff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffdfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 311
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1240: ir 'h%h !== 'hf", ir); end	// Vector No: 310
assert (op === 'hf8) else begin fail = 1; $display("Error 1241: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1242: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1243: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffdfff:1:1:f:f8:0:07ffd:
//------------------------

#2;
word <= 'hffffffffffffdfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 312
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1244: ir 'h%h !== 'hf", ir); end	// Vector No: 311
assert (op === 'hf8) else begin fail = 1; $display("Error 1245: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1246: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffd) else begin fail = 1; $display("Error 1247: addr 'h%h !== 'h07ffd", addr); end
#2;
clk <= 0;

// ffffffffffffbfff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffffbfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 313
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1248: ir 'h%h !== 'hf", ir); end	// Vector No: 312
assert (op === 'hff) else begin fail = 1; $display("Error 1249: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1250: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1251: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffffbfff:0:1:f:ff:0:fbfff:
//------------------------

#2;
word <= 'hffffffffffffbfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 314
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1252: ir 'h%h !== 'hf", ir); end	// Vector No: 313
assert (op === 'hff) else begin fail = 1; $display("Error 1253: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1254: extop 'h%h !== 0", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 1255: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// ffffffffffffbfff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffffbfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 315
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1256: ir 'h%h !== 'hf", ir); end	// Vector No: 314
assert (op === 'hf8) else begin fail = 1; $display("Error 1257: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1258: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1259: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffffbfff:1:1:f:f8:0:07ffb:
//------------------------

#2;
word <= 'hffffffffffffbfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 316
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1260: ir 'h%h !== 'hf", ir); end	// Vector No: 315
assert (op === 'hf8) else begin fail = 1; $display("Error 1261: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1262: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffb) else begin fail = 1; $display("Error 1263: addr 'h%h !== 'h07ffb", addr); end
#2;
clk <= 0;

// ffffffffffff7fff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffff7fff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 317
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1264: ir 'h%h !== 'hf", ir); end	// Vector No: 316
assert (op === 'hff) else begin fail = 1; $display("Error 1265: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1266: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1267: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffff7fff:0:1:f:ff:0:f7fff:
//------------------------

#2;
word <= 'hffffffffffff7fff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 318
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1268: ir 'h%h !== 'hf", ir); end	// Vector No: 317
assert (op === 'hff) else begin fail = 1; $display("Error 1269: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1270: extop 'h%h !== 0", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 1271: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// ffffffffffff7fff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffff7fff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 319
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1272: ir 'h%h !== 'hf", ir); end	// Vector No: 318
assert (op === 'hf8) else begin fail = 1; $display("Error 1273: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1274: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1275: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffff7fff:1:1:f:f8:0:07ff7:
//------------------------

#2;
word <= 'hffffffffffff7fff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 320
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1276: ir 'h%h !== 'hf", ir); end	// Vector No: 319
assert (op === 'hf8) else begin fail = 1; $display("Error 1277: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1278: extop 'h%h !== 0", extop); end
assert (addr === 'h07ff7) else begin fail = 1; $display("Error 1279: addr 'h%h !== 'h07ff7", addr); end
#2;
clk <= 0;

// fffffffffffeffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffeffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 321
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1280: ir 'h%h !== 'hf", ir); end	// Vector No: 320
assert (op === 'hff) else begin fail = 1; $display("Error 1281: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1282: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1283: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffeffff:0:1:f:ff:0:effff:
//------------------------

#2;
word <= 'hfffffffffffeffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 322
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1284: ir 'h%h !== 'hf", ir); end	// Vector No: 321
assert (op === 'hff) else begin fail = 1; $display("Error 1285: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1286: extop 'h%h !== 0", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 1287: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// fffffffffffeffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffeffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 323
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1288: ir 'h%h !== 'hf", ir); end	// Vector No: 322
assert (op === 'hf8) else begin fail = 1; $display("Error 1289: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1290: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1291: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffeffff:1:1:f:f8:0:07fef:
//------------------------

#2;
word <= 'hfffffffffffeffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 324
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1292: ir 'h%h !== 'hf", ir); end	// Vector No: 323
assert (op === 'hf8) else begin fail = 1; $display("Error 1293: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1294: extop 'h%h !== 0", extop); end
assert (addr === 'h07fef) else begin fail = 1; $display("Error 1295: addr 'h%h !== 'h07fef", addr); end
#2;
clk <= 0;

// fffffffffffdffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffdffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 325
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1296: ir 'h%h !== 'hf", ir); end	// Vector No: 324
assert (op === 'hff) else begin fail = 1; $display("Error 1297: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1298: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1299: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffdffff:0:1:f:ff:0:dffff:
//------------------------

#2;
word <= 'hfffffffffffdffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 326
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1300: ir 'h%h !== 'hf", ir); end	// Vector No: 325
assert (op === 'hff) else begin fail = 1; $display("Error 1301: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1302: extop 'h%h !== 0", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 1303: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// fffffffffffdffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffdffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 327
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1304: ir 'h%h !== 'hf", ir); end	// Vector No: 326
assert (op === 'hf8) else begin fail = 1; $display("Error 1305: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1306: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1307: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffdffff:1:1:f:f8:0:07fdf:
//------------------------

#2;
word <= 'hfffffffffffdffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 328
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1308: ir 'h%h !== 'hf", ir); end	// Vector No: 327
assert (op === 'hf8) else begin fail = 1; $display("Error 1309: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1310: extop 'h%h !== 0", extop); end
assert (addr === 'h07fdf) else begin fail = 1; $display("Error 1311: addr 'h%h !== 'h07fdf", addr); end
#2;
clk <= 0;

// fffffffffffbffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffffbffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 329
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1312: ir 'h%h !== 'hf", ir); end	// Vector No: 328
assert (op === 'hff) else begin fail = 1; $display("Error 1313: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1314: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1315: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffffbffff:0:1:f:ff:0:bffff:
//------------------------

#2;
word <= 'hfffffffffffbffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 330
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1316: ir 'h%h !== 'hf", ir); end	// Vector No: 329
assert (op === 'hff) else begin fail = 1; $display("Error 1317: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1318: extop 'h%h !== 0", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 1319: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// fffffffffffbffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffffbffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 331
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1320: ir 'h%h !== 'hf", ir); end	// Vector No: 330
assert (op === 'hf8) else begin fail = 1; $display("Error 1321: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1322: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1323: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffffbffff:1:1:f:f8:0:07fbf:
//------------------------

#2;
word <= 'hfffffffffffbffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 332
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1324: ir 'h%h !== 'hf", ir); end	// Vector No: 331
assert (op === 'hf8) else begin fail = 1; $display("Error 1325: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1326: extop 'h%h !== 0", extop); end
assert (addr === 'h07fbf) else begin fail = 1; $display("Error 1327: addr 'h%h !== 'h07fbf", addr); end
#2;
clk <= 0;

// fffffffffff7ffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffff7ffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 333
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1328: ir 'h%h !== 'hf", ir); end	// Vector No: 332
assert (op === 'hff) else begin fail = 1; $display("Error 1329: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1330: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1331: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffff7ffff:0:1:f:ff:0:7ffff:
//------------------------

#2;
word <= 'hfffffffffff7ffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 334
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1332: ir 'h%h !== 'hf", ir); end	// Vector No: 333
assert (op === 'hff) else begin fail = 1; $display("Error 1333: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1334: extop 'h%h !== 0", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 1335: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// fffffffffff7ffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffff7ffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 335
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1336: ir 'h%h !== 'hf", ir); end	// Vector No: 334
assert (op === 'hf8) else begin fail = 1; $display("Error 1337: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1338: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1339: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffff7ffff:1:1:f:f8:0:07f7f:
//------------------------

#2;
word <= 'hfffffffffff7ffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 336
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1340: ir 'h%h !== 'hf", ir); end	// Vector No: 335
assert (op === 'hf8) else begin fail = 1; $display("Error 1341: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1342: extop 'h%h !== 0", extop); end
assert (addr === 'h07f7f) else begin fail = 1; $display("Error 1343: addr 'h%h !== 'h07f7f", addr); end
#2;
clk <= 0;

// ffffffffffefffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffefffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 337
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1344: ir 'h%h !== 'hf", ir); end	// Vector No: 336
assert (op === 'hff) else begin fail = 1; $display("Error 1345: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1346: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1347: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffefffff:0:1:f:fe:0:fffff:
//------------------------

#2;
word <= 'hffffffffffefffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 338
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1348: ir 'h%h !== 'hf", ir); end	// Vector No: 337
assert (op === 'hfe) else begin fail = 1; $display("Error 1349: op 'h%h !== 'hfe", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1350: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1351: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffefffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffefffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 339
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1352: ir 'h%h !== 'hf", ir); end	// Vector No: 338
assert (op === 'hf8) else begin fail = 1; $display("Error 1353: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1354: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1355: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffefffff:1:1:f:f8:0:07eff:
//------------------------

#2;
word <= 'hffffffffffefffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 340
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1356: ir 'h%h !== 'hf", ir); end	// Vector No: 339
assert (op === 'hf8) else begin fail = 1; $display("Error 1357: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1358: extop 'h%h !== 0", extop); end
assert (addr === 'h07eff) else begin fail = 1; $display("Error 1359: addr 'h%h !== 'h07eff", addr); end
#2;
clk <= 0;

// ffffffffffdfffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffdfffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 341
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1360: ir 'h%h !== 'hf", ir); end	// Vector No: 340
assert (op === 'hff) else begin fail = 1; $display("Error 1361: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1362: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1363: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffdfffff:0:1:f:fd:0:fffff:
//------------------------

#2;
word <= 'hffffffffffdfffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 342
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1364: ir 'h%h !== 'hf", ir); end	// Vector No: 341
assert (op === 'hfd) else begin fail = 1; $display("Error 1365: op 'h%h !== 'hfd", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1366: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1367: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffdfffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffdfffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 343
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1368: ir 'h%h !== 'hf", ir); end	// Vector No: 342
assert (op === 'hf8) else begin fail = 1; $display("Error 1369: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1370: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1371: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffdfffff:1:1:f:f8:0:07dff:
//------------------------

#2;
word <= 'hffffffffffdfffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 344
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1372: ir 'h%h !== 'hf", ir); end	// Vector No: 343
assert (op === 'hf8) else begin fail = 1; $display("Error 1373: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1374: extop 'h%h !== 0", extop); end
assert (addr === 'h07dff) else begin fail = 1; $display("Error 1375: addr 'h%h !== 'h07dff", addr); end
#2;
clk <= 0;

// ffffffffffbfffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffffbfffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 345
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1376: ir 'h%h !== 'hf", ir); end	// Vector No: 344
assert (op === 'hff) else begin fail = 1; $display("Error 1377: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1378: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1379: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffbfffff:0:1:f:fb:0:fffff:
//------------------------

#2;
word <= 'hffffffffffbfffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 346
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1380: ir 'h%h !== 'hf", ir); end	// Vector No: 345
assert (op === 'hfb) else begin fail = 1; $display("Error 1381: op 'h%h !== 'hfb", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1382: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1383: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffffbfffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffffbfffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 347
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1384: ir 'h%h !== 'hf", ir); end	// Vector No: 346
assert (op === 'hf8) else begin fail = 1; $display("Error 1385: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1386: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1387: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffffbfffff:1:1:f:f8:0:07bff:
//------------------------

#2;
word <= 'hffffffffffbfffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 348
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1388: ir 'h%h !== 'hf", ir); end	// Vector No: 347
assert (op === 'hf8) else begin fail = 1; $display("Error 1389: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1390: extop 'h%h !== 0", extop); end
assert (addr === 'h07bff) else begin fail = 1; $display("Error 1391: addr 'h%h !== 'h07bff", addr); end
#2;
clk <= 0;

// ffffffffff7fffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffff7fffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 349
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1392: ir 'h%h !== 'hf", ir); end	// Vector No: 348
assert (op === 'hff) else begin fail = 1; $display("Error 1393: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1394: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1395: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffff7fffff:0:1:f:f7:0:fffff:
//------------------------

#2;
word <= 'hffffffffff7fffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 350
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1396: ir 'h%h !== 'hf", ir); end	// Vector No: 349
assert (op === 'hf7) else begin fail = 1; $display("Error 1397: op 'h%h !== 'hf7", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1398: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1399: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffff7fffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffff7fffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 351
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1400: ir 'h%h !== 'hf", ir); end	// Vector No: 350
assert (op === 'hf8) else begin fail = 1; $display("Error 1401: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1402: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1403: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffff7fffff:1:1:f:f8:0:077ff:
//------------------------

#2;
word <= 'hffffffffff7fffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 352
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1404: ir 'h%h !== 'hf", ir); end	// Vector No: 351
assert (op === 'hf8) else begin fail = 1; $display("Error 1405: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1406: extop 'h%h !== 0", extop); end
assert (addr === 'h077ff) else begin fail = 1; $display("Error 1407: addr 'h%h !== 'h077ff", addr); end
#2;
clk <= 0;

// fffffffffeffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffeffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 353
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1408: ir 'h%h !== 'hf", ir); end	// Vector No: 352
assert (op === 'hff) else begin fail = 1; $display("Error 1409: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1410: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1411: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffeffffff:0:1:f:ef:0:fffff:
//------------------------

#2;
word <= 'hfffffffffeffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 354
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1412: ir 'h%h !== 'hf", ir); end	// Vector No: 353
assert (op === 'hef) else begin fail = 1; $display("Error 1413: op 'h%h !== 'hef", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1414: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1415: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffeffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffeffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 355
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1416: ir 'h%h !== 'hf", ir); end	// Vector No: 354
assert (op === 'hf8) else begin fail = 1; $display("Error 1417: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1418: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1419: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffeffffff:1:1:f:f8:0:06fff:
//------------------------

#2;
word <= 'hfffffffffeffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 356
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1420: ir 'h%h !== 'hf", ir); end	// Vector No: 355
assert (op === 'hf8) else begin fail = 1; $display("Error 1421: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1422: extop 'h%h !== 0", extop); end
assert (addr === 'h06fff) else begin fail = 1; $display("Error 1423: addr 'h%h !== 'h06fff", addr); end
#2;
clk <= 0;

// fffffffffdffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffdffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 357
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1424: ir 'h%h !== 'hf", ir); end	// Vector No: 356
assert (op === 'hff) else begin fail = 1; $display("Error 1425: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1426: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1427: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffdffffff:0:1:f:df:0:fffff:
//------------------------

#2;
word <= 'hfffffffffdffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 358
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1428: ir 'h%h !== 'hf", ir); end	// Vector No: 357
assert (op === 'hdf) else begin fail = 1; $display("Error 1429: op 'h%h !== 'hdf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1430: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1431: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffdffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffdffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 359
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1432: ir 'h%h !== 'hf", ir); end	// Vector No: 358
assert (op === 'hf8) else begin fail = 1; $display("Error 1433: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1434: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1435: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffdffffff:1:1:f:f8:0:05fff:
//------------------------

#2;
word <= 'hfffffffffdffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 360
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1436: ir 'h%h !== 'hf", ir); end	// Vector No: 359
assert (op === 'hf8) else begin fail = 1; $display("Error 1437: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1438: extop 'h%h !== 0", extop); end
assert (addr === 'h05fff) else begin fail = 1; $display("Error 1439: addr 'h%h !== 'h05fff", addr); end
#2;
clk <= 0;

// fffffffffbffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffffbffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 361
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1440: ir 'h%h !== 'hf", ir); end	// Vector No: 360
assert (op === 'hff) else begin fail = 1; $display("Error 1441: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1442: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1443: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffbffffff:0:1:f:bf:0:fffff:
//------------------------

#2;
word <= 'hfffffffffbffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 362
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1444: ir 'h%h !== 'hf", ir); end	// Vector No: 361
assert (op === 'hbf) else begin fail = 1; $display("Error 1445: op 'h%h !== 'hbf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1446: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1447: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffffbffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffffbffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 363
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1448: ir 'h%h !== 'hf", ir); end	// Vector No: 362
assert (op === 'hf8) else begin fail = 1; $display("Error 1449: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1450: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1451: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffffbffffff:1:1:f:f8:0:03fff:
//------------------------

#2;
word <= 'hfffffffffbffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 364
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1452: ir 'h%h !== 'hf", ir); end	// Vector No: 363
assert (op === 'hf8) else begin fail = 1; $display("Error 1453: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1454: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 1455: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fffffffff7ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff7ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 365
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1456: ir 'h%h !== 'hf", ir); end	// Vector No: 364
assert (op === 'hff) else begin fail = 1; $display("Error 1457: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1458: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1459: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff7ffffff:0:1:f:7f:0:fffff:
//------------------------

#2;
word <= 'hfffffffff7ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 366
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1460: ir 'h%h !== 'hf", ir); end	// Vector No: 365
assert (op === 'h7f) else begin fail = 1; $display("Error 1461: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1462: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1463: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff7ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff7ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 367
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1464: ir 'h%h !== 'hf", ir); end	// Vector No: 366
assert (op === 'hf8) else begin fail = 1; $display("Error 1465: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1466: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1467: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff7ffffff:1:1:f:f0:0:07fff:
//------------------------

#2;
word <= 'hfffffffff7ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 368
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1468: ir 'h%h !== 'hf", ir); end	// Vector No: 367
assert (op === 'hf0) else begin fail = 1; $display("Error 1469: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1470: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1471: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffefffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffefffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 369
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1472: ir 'h%h !== 'hf", ir); end	// Vector No: 368
assert (op === 'hff) else begin fail = 1; $display("Error 1473: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1474: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1475: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffefffffff:0:1:e:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffefffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 370
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 1476: ir 'h%h !== 'he", ir); end	// Vector No: 369
assert (op === 'hff) else begin fail = 1; $display("Error 1477: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1478: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1479: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffefffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffefffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 371
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1480: ir 'h%h !== 'hf", ir); end	// Vector No: 370
assert (op === 'hf8) else begin fail = 1; $display("Error 1481: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1482: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1483: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffefffffff:1:1:f:e8:0:07fff:
//------------------------

#2;
word <= 'hffffffffefffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 372
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1484: ir 'h%h !== 'hf", ir); end	// Vector No: 371
assert (op === 'he8) else begin fail = 1; $display("Error 1485: op 'h%h !== 'he8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1486: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1487: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffdfffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffdfffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 373
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1488: ir 'h%h !== 'hf", ir); end	// Vector No: 372
assert (op === 'hff) else begin fail = 1; $display("Error 1489: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1490: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1491: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffdfffffff:0:1:d:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffdfffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 374
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 1492: ir 'h%h !== 'hd", ir); end	// Vector No: 373
assert (op === 'hff) else begin fail = 1; $display("Error 1493: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1494: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1495: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffdfffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffdfffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 375
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1496: ir 'h%h !== 'hf", ir); end	// Vector No: 374
assert (op === 'hf8) else begin fail = 1; $display("Error 1497: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1498: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1499: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffdfffffff:1:1:f:d8:0:07fff:
//------------------------

#2;
word <= 'hffffffffdfffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 376
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1500: ir 'h%h !== 'hf", ir); end	// Vector No: 375
assert (op === 'hd8) else begin fail = 1; $display("Error 1501: op 'h%h !== 'hd8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1502: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1503: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffbfffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffbfffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 377
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1504: ir 'h%h !== 'hf", ir); end	// Vector No: 376
assert (op === 'hff) else begin fail = 1; $display("Error 1505: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1506: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1507: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffbfffffff:0:1:b:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffbfffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 378
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 1508: ir 'h%h !== 'hb", ir); end	// Vector No: 377
assert (op === 'hff) else begin fail = 1; $display("Error 1509: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1510: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1511: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffbfffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffbfffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 379
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1512: ir 'h%h !== 'hf", ir); end	// Vector No: 378
assert (op === 'hf8) else begin fail = 1; $display("Error 1513: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1514: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1515: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffbfffffff:1:1:f:b8:0:07fff:
//------------------------

#2;
word <= 'hffffffffbfffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 380
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1516: ir 'h%h !== 'hf", ir); end	// Vector No: 379
assert (op === 'hb8) else begin fail = 1; $display("Error 1517: op 'h%h !== 'hb8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1518: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1519: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffff7fffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffff7fffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 381
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1520: ir 'h%h !== 'hf", ir); end	// Vector No: 380
assert (op === 'hff) else begin fail = 1; $display("Error 1521: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1522: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1523: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffff7fffffff:0:1:7:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffff7fffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 382
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 1524: ir 'h%h !== 'h7", ir); end	// Vector No: 381
assert (op === 'hff) else begin fail = 1; $display("Error 1525: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1526: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1527: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffff7fffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffff7fffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 383
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1528: ir 'h%h !== 'hf", ir); end	// Vector No: 382
assert (op === 'hf8) else begin fail = 1; $display("Error 1529: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1530: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1531: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffff7fffffff:1:1:f:7f:0:07fff:
//------------------------

#2;
word <= 'hffffffff7fffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 384
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1532: ir 'h%h !== 'hf", ir); end	// Vector No: 383
assert (op === 'h7f) else begin fail = 1; $display("Error 1533: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1534: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1535: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffeffffffff:0:0:f:ff:0:ffffe:
//------------------------

#2;
word <= 'hfffffffeffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 385
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1536: ir 'h%h !== 'hf", ir); end	// Vector No: 384
assert (op === 'hff) else begin fail = 1; $display("Error 1537: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1538: extop 'h%h !== 0", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 1539: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// fffffffeffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffeffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 386
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1540: ir 'h%h !== 'hf", ir); end	// Vector No: 385
assert (op === 'hff) else begin fail = 1; $display("Error 1541: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1542: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1543: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffeffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffeffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 387
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1544: ir 'h%h !== 'hf", ir); end	// Vector No: 386
assert (op === 'hf8) else begin fail = 1; $display("Error 1545: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1546: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1547: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffeffffffff:1:1:e:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffeffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 388
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 1548: ir 'h%h !== 'he", ir); end	// Vector No: 387
assert (op === 'hf8) else begin fail = 1; $display("Error 1549: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1550: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1551: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffdffffffff:0:0:f:ff:0:ffffd:
//------------------------

#2;
word <= 'hfffffffdffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 389
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1552: ir 'h%h !== 'hf", ir); end	// Vector No: 388
assert (op === 'hff) else begin fail = 1; $display("Error 1553: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1554: extop 'h%h !== 0", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 1555: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// fffffffdffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffdffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 390
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1556: ir 'h%h !== 'hf", ir); end	// Vector No: 389
assert (op === 'hff) else begin fail = 1; $display("Error 1557: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1558: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1559: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffdffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffdffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 391
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1560: ir 'h%h !== 'hf", ir); end	// Vector No: 390
assert (op === 'hf8) else begin fail = 1; $display("Error 1561: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1562: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1563: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffdffffffff:1:1:d:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffdffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 392
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 1564: ir 'h%h !== 'hd", ir); end	// Vector No: 391
assert (op === 'hf8) else begin fail = 1; $display("Error 1565: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1566: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1567: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffbffffffff:0:0:f:ff:0:ffffb:
//------------------------

#2;
word <= 'hfffffffbffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 393
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1568: ir 'h%h !== 'hf", ir); end	// Vector No: 392
assert (op === 'hff) else begin fail = 1; $display("Error 1569: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1570: extop 'h%h !== 0", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 1571: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// fffffffbffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffbffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 394
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1572: ir 'h%h !== 'hf", ir); end	// Vector No: 393
assert (op === 'hff) else begin fail = 1; $display("Error 1573: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1574: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1575: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffbffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffbffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 395
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1576: ir 'h%h !== 'hf", ir); end	// Vector No: 394
assert (op === 'hf8) else begin fail = 1; $display("Error 1577: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1578: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1579: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffbffffffff:1:1:b:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffbffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 396
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 1580: ir 'h%h !== 'hb", ir); end	// Vector No: 395
assert (op === 'hf8) else begin fail = 1; $display("Error 1581: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1582: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1583: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffff7ffffffff:0:0:f:ff:0:ffff7:
//------------------------

#2;
word <= 'hfffffff7ffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 397
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1584: ir 'h%h !== 'hf", ir); end	// Vector No: 396
assert (op === 'hff) else begin fail = 1; $display("Error 1585: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1586: extop 'h%h !== 0", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 1587: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// fffffff7ffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffff7ffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 398
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1588: ir 'h%h !== 'hf", ir); end	// Vector No: 397
assert (op === 'hff) else begin fail = 1; $display("Error 1589: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1590: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1591: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffff7ffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffff7ffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 399
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1592: ir 'h%h !== 'hf", ir); end	// Vector No: 398
assert (op === 'hf8) else begin fail = 1; $display("Error 1593: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1594: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1595: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffff7ffffffff:1:1:7:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffff7ffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 400
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 1596: ir 'h%h !== 'h7", ir); end	// Vector No: 399
assert (op === 'hf8) else begin fail = 1; $display("Error 1597: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1598: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1599: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffefffffffff:0:0:f:ff:0:fffef:
//------------------------

#2;
word <= 'hffffffefffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 401
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1600: ir 'h%h !== 'hf", ir); end	// Vector No: 400
assert (op === 'hff) else begin fail = 1; $display("Error 1601: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1602: extop 'h%h !== 0", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 1603: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// ffffffefffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffefffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 402
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1604: ir 'h%h !== 'hf", ir); end	// Vector No: 401
assert (op === 'hff) else begin fail = 1; $display("Error 1605: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1606: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1607: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffefffffffff:1:0:f:f8:0:07ffe:
//------------------------

#2;
word <= 'hffffffefffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 403
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1608: ir 'h%h !== 'hf", ir); end	// Vector No: 402
assert (op === 'hf8) else begin fail = 1; $display("Error 1609: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1610: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffe) else begin fail = 1; $display("Error 1611: addr 'h%h !== 'h07ffe", addr); end
#2;
clk <= 0;

// ffffffefffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffefffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 404
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1612: ir 'h%h !== 'hf", ir); end	// Vector No: 403
assert (op === 'hf8) else begin fail = 1; $display("Error 1613: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1614: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1615: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffdfffffffff:0:0:f:ff:0:fffdf:
//------------------------

#2;
word <= 'hffffffdfffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 405
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1616: ir 'h%h !== 'hf", ir); end	// Vector No: 404
assert (op === 'hff) else begin fail = 1; $display("Error 1617: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1618: extop 'h%h !== 0", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 1619: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// ffffffdfffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffdfffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 406
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1620: ir 'h%h !== 'hf", ir); end	// Vector No: 405
assert (op === 'hff) else begin fail = 1; $display("Error 1621: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1622: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1623: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffdfffffffff:1:0:f:f8:0:07ffd:
//------------------------

#2;
word <= 'hffffffdfffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 407
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1624: ir 'h%h !== 'hf", ir); end	// Vector No: 406
assert (op === 'hf8) else begin fail = 1; $display("Error 1625: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1626: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffd) else begin fail = 1; $display("Error 1627: addr 'h%h !== 'h07ffd", addr); end
#2;
clk <= 0;

// ffffffdfffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffdfffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 408
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1628: ir 'h%h !== 'hf", ir); end	// Vector No: 407
assert (op === 'hf8) else begin fail = 1; $display("Error 1629: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1630: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1631: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffbfffffffff:0:0:f:ff:0:fffbf:
//------------------------

#2;
word <= 'hffffffbfffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 409
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1632: ir 'h%h !== 'hf", ir); end	// Vector No: 408
assert (op === 'hff) else begin fail = 1; $display("Error 1633: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1634: extop 'h%h !== 0", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 1635: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// ffffffbfffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffbfffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 410
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1636: ir 'h%h !== 'hf", ir); end	// Vector No: 409
assert (op === 'hff) else begin fail = 1; $display("Error 1637: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1638: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1639: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffbfffffffff:1:0:f:f8:0:07ffb:
//------------------------

#2;
word <= 'hffffffbfffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 411
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1640: ir 'h%h !== 'hf", ir); end	// Vector No: 410
assert (op === 'hf8) else begin fail = 1; $display("Error 1641: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1642: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffb) else begin fail = 1; $display("Error 1643: addr 'h%h !== 'h07ffb", addr); end
#2;
clk <= 0;

// ffffffbfffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffbfffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 412
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1644: ir 'h%h !== 'hf", ir); end	// Vector No: 411
assert (op === 'hf8) else begin fail = 1; $display("Error 1645: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1646: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1647: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffff7fffffffff:0:0:f:ff:0:fff7f:
//------------------------

#2;
word <= 'hffffff7fffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 413
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1648: ir 'h%h !== 'hf", ir); end	// Vector No: 412
assert (op === 'hff) else begin fail = 1; $display("Error 1649: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1650: extop 'h%h !== 0", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 1651: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// ffffff7fffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffff7fffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 414
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1652: ir 'h%h !== 'hf", ir); end	// Vector No: 413
assert (op === 'hff) else begin fail = 1; $display("Error 1653: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1654: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1655: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffff7fffffffff:1:0:f:f8:0:07ff7:
//------------------------

#2;
word <= 'hffffff7fffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 415
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1656: ir 'h%h !== 'hf", ir); end	// Vector No: 414
assert (op === 'hf8) else begin fail = 1; $display("Error 1657: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1658: extop 'h%h !== 0", extop); end
assert (addr === 'h07ff7) else begin fail = 1; $display("Error 1659: addr 'h%h !== 'h07ff7", addr); end
#2;
clk <= 0;

// ffffff7fffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffff7fffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 416
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1660: ir 'h%h !== 'hf", ir); end	// Vector No: 415
assert (op === 'hf8) else begin fail = 1; $display("Error 1661: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1662: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1663: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffeffffffffff:0:0:f:ff:0:ffeff:
//------------------------

#2;
word <= 'hfffffeffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 417
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1664: ir 'h%h !== 'hf", ir); end	// Vector No: 416
assert (op === 'hff) else begin fail = 1; $display("Error 1665: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1666: extop 'h%h !== 0", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 1667: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// fffffeffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffeffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 418
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1668: ir 'h%h !== 'hf", ir); end	// Vector No: 417
assert (op === 'hff) else begin fail = 1; $display("Error 1669: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1670: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1671: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffeffffffffff:1:0:f:f8:0:07fef:
//------------------------

#2;
word <= 'hfffffeffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 419
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1672: ir 'h%h !== 'hf", ir); end	// Vector No: 418
assert (op === 'hf8) else begin fail = 1; $display("Error 1673: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1674: extop 'h%h !== 0", extop); end
assert (addr === 'h07fef) else begin fail = 1; $display("Error 1675: addr 'h%h !== 'h07fef", addr); end
#2;
clk <= 0;

// fffffeffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffeffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 420
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1676: ir 'h%h !== 'hf", ir); end	// Vector No: 419
assert (op === 'hf8) else begin fail = 1; $display("Error 1677: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1678: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1679: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffdffffffffff:0:0:f:ff:0:ffdff:
//------------------------

#2;
word <= 'hfffffdffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 421
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1680: ir 'h%h !== 'hf", ir); end	// Vector No: 420
assert (op === 'hff) else begin fail = 1; $display("Error 1681: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1682: extop 'h%h !== 0", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 1683: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// fffffdffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffdffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 422
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1684: ir 'h%h !== 'hf", ir); end	// Vector No: 421
assert (op === 'hff) else begin fail = 1; $display("Error 1685: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1686: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1687: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffdffffffffff:1:0:f:f8:0:07fdf:
//------------------------

#2;
word <= 'hfffffdffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 423
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1688: ir 'h%h !== 'hf", ir); end	// Vector No: 422
assert (op === 'hf8) else begin fail = 1; $display("Error 1689: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1690: extop 'h%h !== 0", extop); end
assert (addr === 'h07fdf) else begin fail = 1; $display("Error 1691: addr 'h%h !== 'h07fdf", addr); end
#2;
clk <= 0;

// fffffdffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffdffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 424
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1692: ir 'h%h !== 'hf", ir); end	// Vector No: 423
assert (op === 'hf8) else begin fail = 1; $display("Error 1693: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1694: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1695: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffbffffffffff:0:0:f:ff:0:ffbff:
//------------------------

#2;
word <= 'hfffffbffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 425
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1696: ir 'h%h !== 'hf", ir); end	// Vector No: 424
assert (op === 'hff) else begin fail = 1; $display("Error 1697: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1698: extop 'h%h !== 0", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 1699: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// fffffbffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffbffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 426
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1700: ir 'h%h !== 'hf", ir); end	// Vector No: 425
assert (op === 'hff) else begin fail = 1; $display("Error 1701: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1702: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1703: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffbffffffffff:1:0:f:f8:0:07fbf:
//------------------------

#2;
word <= 'hfffffbffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 427
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1704: ir 'h%h !== 'hf", ir); end	// Vector No: 426
assert (op === 'hf8) else begin fail = 1; $display("Error 1705: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1706: extop 'h%h !== 0", extop); end
assert (addr === 'h07fbf) else begin fail = 1; $display("Error 1707: addr 'h%h !== 'h07fbf", addr); end
#2;
clk <= 0;

// fffffbffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffbffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 428
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1708: ir 'h%h !== 'hf", ir); end	// Vector No: 427
assert (op === 'hf8) else begin fail = 1; $display("Error 1709: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1710: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1711: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffff7ffffffffff:0:0:f:ff:0:ff7ff:
//------------------------

#2;
word <= 'hfffff7ffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 429
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1712: ir 'h%h !== 'hf", ir); end	// Vector No: 428
assert (op === 'hff) else begin fail = 1; $display("Error 1713: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1714: extop 'h%h !== 0", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 1715: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// fffff7ffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffff7ffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 430
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1716: ir 'h%h !== 'hf", ir); end	// Vector No: 429
assert (op === 'hff) else begin fail = 1; $display("Error 1717: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1718: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1719: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffff7ffffffffff:1:0:f:f8:0:07f7f:
//------------------------

#2;
word <= 'hfffff7ffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 431
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1720: ir 'h%h !== 'hf", ir); end	// Vector No: 430
assert (op === 'hf8) else begin fail = 1; $display("Error 1721: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1722: extop 'h%h !== 0", extop); end
assert (addr === 'h07f7f) else begin fail = 1; $display("Error 1723: addr 'h%h !== 'h07f7f", addr); end
#2;
clk <= 0;

// fffff7ffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffff7ffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 432
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1724: ir 'h%h !== 'hf", ir); end	// Vector No: 431
assert (op === 'hf8) else begin fail = 1; $display("Error 1725: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1726: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1727: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffefffffffffff:0:0:f:ff:0:fefff:
//------------------------

#2;
word <= 'hffffefffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 433
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1728: ir 'h%h !== 'hf", ir); end	// Vector No: 432
assert (op === 'hff) else begin fail = 1; $display("Error 1729: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1730: extop 'h%h !== 0", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 1731: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// ffffefffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffefffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 434
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1732: ir 'h%h !== 'hf", ir); end	// Vector No: 433
assert (op === 'hff) else begin fail = 1; $display("Error 1733: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1734: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1735: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffefffffffffff:1:0:f:f8:0:07eff:
//------------------------

#2;
word <= 'hffffefffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 435
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1736: ir 'h%h !== 'hf", ir); end	// Vector No: 434
assert (op === 'hf8) else begin fail = 1; $display("Error 1737: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1738: extop 'h%h !== 0", extop); end
assert (addr === 'h07eff) else begin fail = 1; $display("Error 1739: addr 'h%h !== 'h07eff", addr); end
#2;
clk <= 0;

// ffffefffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffefffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 436
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1740: ir 'h%h !== 'hf", ir); end	// Vector No: 435
assert (op === 'hf8) else begin fail = 1; $display("Error 1741: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1742: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1743: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffdfffffffffff:0:0:f:ff:0:fdfff:
//------------------------

#2;
word <= 'hffffdfffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 437
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1744: ir 'h%h !== 'hf", ir); end	// Vector No: 436
assert (op === 'hff) else begin fail = 1; $display("Error 1745: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1746: extop 'h%h !== 0", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 1747: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// ffffdfffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffdfffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 438
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1748: ir 'h%h !== 'hf", ir); end	// Vector No: 437
assert (op === 'hff) else begin fail = 1; $display("Error 1749: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1750: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1751: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffdfffffffffff:1:0:f:f8:0:07dff:
//------------------------

#2;
word <= 'hffffdfffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 439
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1752: ir 'h%h !== 'hf", ir); end	// Vector No: 438
assert (op === 'hf8) else begin fail = 1; $display("Error 1753: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1754: extop 'h%h !== 0", extop); end
assert (addr === 'h07dff) else begin fail = 1; $display("Error 1755: addr 'h%h !== 'h07dff", addr); end
#2;
clk <= 0;

// ffffdfffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffdfffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 440
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1756: ir 'h%h !== 'hf", ir); end	// Vector No: 439
assert (op === 'hf8) else begin fail = 1; $display("Error 1757: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1758: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1759: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffbfffffffffff:0:0:f:ff:0:fbfff:
//------------------------

#2;
word <= 'hffffbfffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 441
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1760: ir 'h%h !== 'hf", ir); end	// Vector No: 440
assert (op === 'hff) else begin fail = 1; $display("Error 1761: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1762: extop 'h%h !== 0", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 1763: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// ffffbfffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffbfffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 442
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1764: ir 'h%h !== 'hf", ir); end	// Vector No: 441
assert (op === 'hff) else begin fail = 1; $display("Error 1765: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1766: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1767: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffbfffffffffff:1:0:f:f8:0:07bff:
//------------------------

#2;
word <= 'hffffbfffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 443
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1768: ir 'h%h !== 'hf", ir); end	// Vector No: 442
assert (op === 'hf8) else begin fail = 1; $display("Error 1769: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1770: extop 'h%h !== 0", extop); end
assert (addr === 'h07bff) else begin fail = 1; $display("Error 1771: addr 'h%h !== 'h07bff", addr); end
#2;
clk <= 0;

// ffffbfffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffbfffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 444
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1772: ir 'h%h !== 'hf", ir); end	// Vector No: 443
assert (op === 'hf8) else begin fail = 1; $display("Error 1773: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1774: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1775: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffff7fffffffffff:0:0:f:ff:0:f7fff:
//------------------------

#2;
word <= 'hffff7fffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 445
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1776: ir 'h%h !== 'hf", ir); end	// Vector No: 444
assert (op === 'hff) else begin fail = 1; $display("Error 1777: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1778: extop 'h%h !== 0", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 1779: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// ffff7fffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffff7fffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 446
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1780: ir 'h%h !== 'hf", ir); end	// Vector No: 445
assert (op === 'hff) else begin fail = 1; $display("Error 1781: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1782: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1783: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffff7fffffffffff:1:0:f:f8:0:077ff:
//------------------------

#2;
word <= 'hffff7fffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 447
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1784: ir 'h%h !== 'hf", ir); end	// Vector No: 446
assert (op === 'hf8) else begin fail = 1; $display("Error 1785: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1786: extop 'h%h !== 0", extop); end
assert (addr === 'h077ff) else begin fail = 1; $display("Error 1787: addr 'h%h !== 'h077ff", addr); end
#2;
clk <= 0;

// ffff7fffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffff7fffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 448
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1788: ir 'h%h !== 'hf", ir); end	// Vector No: 447
assert (op === 'hf8) else begin fail = 1; $display("Error 1789: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1790: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1791: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffeffffffffffff:0:0:f:ff:0:effff:
//------------------------

#2;
word <= 'hfffeffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 449
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1792: ir 'h%h !== 'hf", ir); end	// Vector No: 448
assert (op === 'hff) else begin fail = 1; $display("Error 1793: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1794: extop 'h%h !== 0", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 1795: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// fffeffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffeffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 450
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1796: ir 'h%h !== 'hf", ir); end	// Vector No: 449
assert (op === 'hff) else begin fail = 1; $display("Error 1797: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1798: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1799: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffeffffffffffff:1:0:f:f8:0:06fff:
//------------------------

#2;
word <= 'hfffeffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 451
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1800: ir 'h%h !== 'hf", ir); end	// Vector No: 450
assert (op === 'hf8) else begin fail = 1; $display("Error 1801: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1802: extop 'h%h !== 0", extop); end
assert (addr === 'h06fff) else begin fail = 1; $display("Error 1803: addr 'h%h !== 'h06fff", addr); end
#2;
clk <= 0;

// fffeffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffeffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 452
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1804: ir 'h%h !== 'hf", ir); end	// Vector No: 451
assert (op === 'hf8) else begin fail = 1; $display("Error 1805: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1806: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1807: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffdffffffffffff:0:0:f:ff:0:dffff:
//------------------------

#2;
word <= 'hfffdffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 453
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1808: ir 'h%h !== 'hf", ir); end	// Vector No: 452
assert (op === 'hff) else begin fail = 1; $display("Error 1809: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1810: extop 'h%h !== 0", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 1811: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// fffdffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffdffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 454
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1812: ir 'h%h !== 'hf", ir); end	// Vector No: 453
assert (op === 'hff) else begin fail = 1; $display("Error 1813: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1814: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1815: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffdffffffffffff:1:0:f:f8:0:05fff:
//------------------------

#2;
word <= 'hfffdffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 455
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1816: ir 'h%h !== 'hf", ir); end	// Vector No: 454
assert (op === 'hf8) else begin fail = 1; $display("Error 1817: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1818: extop 'h%h !== 0", extop); end
assert (addr === 'h05fff) else begin fail = 1; $display("Error 1819: addr 'h%h !== 'h05fff", addr); end
#2;
clk <= 0;

// fffdffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffdffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 456
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1820: ir 'h%h !== 'hf", ir); end	// Vector No: 455
assert (op === 'hf8) else begin fail = 1; $display("Error 1821: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1822: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1823: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffbffffffffffff:0:0:f:ff:0:bffff:
//------------------------

#2;
word <= 'hfffbffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 457
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1824: ir 'h%h !== 'hf", ir); end	// Vector No: 456
assert (op === 'hff) else begin fail = 1; $display("Error 1825: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1826: extop 'h%h !== 0", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 1827: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// fffbffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffbffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 458
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1828: ir 'h%h !== 'hf", ir); end	// Vector No: 457
assert (op === 'hff) else begin fail = 1; $display("Error 1829: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1830: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1831: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffbffffffffffff:1:0:f:f8:0:03fff:
//------------------------

#2;
word <= 'hfffbffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 459
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1832: ir 'h%h !== 'hf", ir); end	// Vector No: 458
assert (op === 'hf8) else begin fail = 1; $display("Error 1833: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1834: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 1835: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fffbffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffbffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 460
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1836: ir 'h%h !== 'hf", ir); end	// Vector No: 459
assert (op === 'hf8) else begin fail = 1; $display("Error 1837: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1838: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1839: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fff7ffffffffffff:0:0:f:ff:0:7ffff:
//------------------------

#2;
word <= 'hfff7ffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 461
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1840: ir 'h%h !== 'hf", ir); end	// Vector No: 460
assert (op === 'hff) else begin fail = 1; $display("Error 1841: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1842: extop 'h%h !== 0", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 1843: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// fff7ffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfff7ffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 462
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1844: ir 'h%h !== 'hf", ir); end	// Vector No: 461
assert (op === 'hff) else begin fail = 1; $display("Error 1845: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1846: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1847: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fff7ffffffffffff:1:0:f:f0:0:07fff:
//------------------------

#2;
word <= 'hfff7ffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 463
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1848: ir 'h%h !== 'hf", ir); end	// Vector No: 462
assert (op === 'hf0) else begin fail = 1; $display("Error 1849: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1850: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1851: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fff7ffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfff7ffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 464
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1852: ir 'h%h !== 'hf", ir); end	// Vector No: 463
assert (op === 'hf8) else begin fail = 1; $display("Error 1853: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1854: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1855: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffefffffffffffff:0:0:f:fe:0:fffff:
//------------------------

#2;
word <= 'hffefffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 465
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1856: ir 'h%h !== 'hf", ir); end	// Vector No: 464
assert (op === 'hfe) else begin fail = 1; $display("Error 1857: op 'h%h !== 'hfe", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1858: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1859: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffefffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffefffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 466
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1860: ir 'h%h !== 'hf", ir); end	// Vector No: 465
assert (op === 'hff) else begin fail = 1; $display("Error 1861: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1862: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1863: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffefffffffffffff:1:0:f:e8:0:07fff:
//------------------------

#2;
word <= 'hffefffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 467
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1864: ir 'h%h !== 'hf", ir); end	// Vector No: 466
assert (op === 'he8) else begin fail = 1; $display("Error 1865: op 'h%h !== 'he8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1866: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1867: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffefffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffefffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 468
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1868: ir 'h%h !== 'hf", ir); end	// Vector No: 467
assert (op === 'hf8) else begin fail = 1; $display("Error 1869: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1870: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1871: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffdfffffffffffff:0:0:f:fd:0:fffff:
//------------------------

#2;
word <= 'hffdfffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 469
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1872: ir 'h%h !== 'hf", ir); end	// Vector No: 468
assert (op === 'hfd) else begin fail = 1; $display("Error 1873: op 'h%h !== 'hfd", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1874: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1875: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffdfffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffdfffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 470
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1876: ir 'h%h !== 'hf", ir); end	// Vector No: 469
assert (op === 'hff) else begin fail = 1; $display("Error 1877: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1878: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1879: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffdfffffffffffff:1:0:f:d8:0:07fff:
//------------------------

#2;
word <= 'hffdfffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 471
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1880: ir 'h%h !== 'hf", ir); end	// Vector No: 470
assert (op === 'hd8) else begin fail = 1; $display("Error 1881: op 'h%h !== 'hd8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1882: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1883: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffdfffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffdfffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 472
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1884: ir 'h%h !== 'hf", ir); end	// Vector No: 471
assert (op === 'hf8) else begin fail = 1; $display("Error 1885: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1886: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1887: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffbfffffffffffff:0:0:f:fb:0:fffff:
//------------------------

#2;
word <= 'hffbfffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 473
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1888: ir 'h%h !== 'hf", ir); end	// Vector No: 472
assert (op === 'hfb) else begin fail = 1; $display("Error 1889: op 'h%h !== 'hfb", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1890: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1891: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffbfffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffbfffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 474
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1892: ir 'h%h !== 'hf", ir); end	// Vector No: 473
assert (op === 'hff) else begin fail = 1; $display("Error 1893: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1894: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1895: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffbfffffffffffff:1:0:f:b8:0:07fff:
//------------------------

#2;
word <= 'hffbfffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 475
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1896: ir 'h%h !== 'hf", ir); end	// Vector No: 474
assert (op === 'hb8) else begin fail = 1; $display("Error 1897: op 'h%h !== 'hb8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1898: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1899: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffbfffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffbfffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 476
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1900: ir 'h%h !== 'hf", ir); end	// Vector No: 475
assert (op === 'hf8) else begin fail = 1; $display("Error 1901: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1902: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1903: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ff7fffffffffffff:0:0:f:f7:0:fffff:
//------------------------

#2;
word <= 'hff7fffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 477
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1904: ir 'h%h !== 'hf", ir); end	// Vector No: 476
assert (op === 'hf7) else begin fail = 1; $display("Error 1905: op 'h%h !== 'hf7", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1906: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1907: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ff7fffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hff7fffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 478
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1908: ir 'h%h !== 'hf", ir); end	// Vector No: 477
assert (op === 'hff) else begin fail = 1; $display("Error 1909: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1910: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1911: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ff7fffffffffffff:1:0:f:7f:0:07fff:
//------------------------

#2;
word <= 'hff7fffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 479
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1912: ir 'h%h !== 'hf", ir); end	// Vector No: 478
assert (op === 'h7f) else begin fail = 1; $display("Error 1913: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1914: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1915: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ff7fffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hff7fffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 480
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1916: ir 'h%h !== 'hf", ir); end	// Vector No: 479
assert (op === 'hf8) else begin fail = 1; $display("Error 1917: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1918: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1919: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// feffffffffffffff:0:0:f:ef:0:fffff:
//------------------------

#2;
word <= 'hfeffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 481
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1920: ir 'h%h !== 'hf", ir); end	// Vector No: 480
assert (op === 'hef) else begin fail = 1; $display("Error 1921: op 'h%h !== 'hef", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1922: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1923: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// feffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfeffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 482
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1924: ir 'h%h !== 'hf", ir); end	// Vector No: 481
assert (op === 'hff) else begin fail = 1; $display("Error 1925: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1926: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1927: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// feffffffffffffff:1:0:e:f8:0:07fff:
//------------------------

#2;
word <= 'hfeffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 483
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 1928: ir 'h%h !== 'he", ir); end	// Vector No: 482
assert (op === 'hf8) else begin fail = 1; $display("Error 1929: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1930: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1931: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// feffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfeffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 484
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1932: ir 'h%h !== 'hf", ir); end	// Vector No: 483
assert (op === 'hf8) else begin fail = 1; $display("Error 1933: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1934: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1935: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fdffffffffffffff:0:0:f:df:0:fffff:
//------------------------

#2;
word <= 'hfdffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 485
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1936: ir 'h%h !== 'hf", ir); end	// Vector No: 484
assert (op === 'hdf) else begin fail = 1; $display("Error 1937: op 'h%h !== 'hdf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1938: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1939: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fdffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfdffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 486
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1940: ir 'h%h !== 'hf", ir); end	// Vector No: 485
assert (op === 'hff) else begin fail = 1; $display("Error 1941: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1942: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1943: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fdffffffffffffff:1:0:d:f8:0:07fff:
//------------------------

#2;
word <= 'hfdffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 487
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 1944: ir 'h%h !== 'hd", ir); end	// Vector No: 486
assert (op === 'hf8) else begin fail = 1; $display("Error 1945: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1946: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1947: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fdffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfdffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 488
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1948: ir 'h%h !== 'hf", ir); end	// Vector No: 487
assert (op === 'hf8) else begin fail = 1; $display("Error 1949: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1950: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1951: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fbffffffffffffff:0:0:f:bf:0:fffff:
//------------------------

#2;
word <= 'hfbffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 489
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1952: ir 'h%h !== 'hf", ir); end	// Vector No: 488
assert (op === 'hbf) else begin fail = 1; $display("Error 1953: op 'h%h !== 'hbf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1954: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1955: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fbffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfbffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 490
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1956: ir 'h%h !== 'hf", ir); end	// Vector No: 489
assert (op === 'hff) else begin fail = 1; $display("Error 1957: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1958: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1959: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fbffffffffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hfbffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 491
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 1960: ir 'h%h !== 'hb", ir); end	// Vector No: 490
assert (op === 'hf8) else begin fail = 1; $display("Error 1961: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1962: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1963: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fbffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfbffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 492
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1964: ir 'h%h !== 'hf", ir); end	// Vector No: 491
assert (op === 'hf8) else begin fail = 1; $display("Error 1965: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1966: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1967: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f7ffffffffffffff:0:0:f:7f:0:fffff:
//------------------------

#2;
word <= 'hf7ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 493
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1968: ir 'h%h !== 'hf", ir); end	// Vector No: 492
assert (op === 'h7f) else begin fail = 1; $display("Error 1969: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1970: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1971: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f7ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf7ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 494
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1972: ir 'h%h !== 'hf", ir); end	// Vector No: 493
assert (op === 'hff) else begin fail = 1; $display("Error 1973: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1974: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1975: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f7ffffffffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf7ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 495
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1976: ir 'h%h !== 'hf", ir); end	// Vector No: 494
assert (op === 'hf8) else begin fail = 1; $display("Error 1977: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1978: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1979: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f7ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf7ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 496
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1980: ir 'h%h !== 'hf", ir); end	// Vector No: 495
assert (op === 'hf8) else begin fail = 1; $display("Error 1981: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1982: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1983: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// efffffffffffffff:0:0:e:ff:0:fffff:
//------------------------

#2;
word <= 'hefffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 497
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 1984: ir 'h%h !== 'he", ir); end	// Vector No: 496
assert (op === 'hff) else begin fail = 1; $display("Error 1985: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1986: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1987: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// efffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hefffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 498
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1988: ir 'h%h !== 'hf", ir); end	// Vector No: 497
assert (op === 'hff) else begin fail = 1; $display("Error 1989: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1990: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 1991: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// efffffffffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hefffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 499
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1992: ir 'h%h !== 'hf", ir); end	// Vector No: 498
assert (op === 'hf8) else begin fail = 1; $display("Error 1993: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1994: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1995: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// efffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hefffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 500
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 1996: ir 'h%h !== 'hf", ir); end	// Vector No: 499
assert (op === 'hf8) else begin fail = 1; $display("Error 1997: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 1998: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 1999: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// dfffffffffffffff:0:0:d:ff:0:fffff:
//------------------------

#2;
word <= 'hdfffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 501
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 2000: ir 'h%h !== 'hd", ir); end	// Vector No: 500
assert (op === 'hff) else begin fail = 1; $display("Error 2001: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2002: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2003: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// dfffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hdfffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 502
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2004: ir 'h%h !== 'hf", ir); end	// Vector No: 501
assert (op === 'hff) else begin fail = 1; $display("Error 2005: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2006: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2007: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// dfffffffffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hdfffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 503
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2008: ir 'h%h !== 'hf", ir); end	// Vector No: 502
assert (op === 'hf8) else begin fail = 1; $display("Error 2009: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2010: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2011: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// dfffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hdfffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 504
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2012: ir 'h%h !== 'hf", ir); end	// Vector No: 503
assert (op === 'hf8) else begin fail = 1; $display("Error 2013: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2014: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2015: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// bfffffffffffffff:0:0:b:ff:0:fffff:
//------------------------

#2;
word <= 'hbfffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 505
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 2016: ir 'h%h !== 'hb", ir); end	// Vector No: 504
assert (op === 'hff) else begin fail = 1; $display("Error 2017: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2018: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2019: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// bfffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hbfffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 506
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2020: ir 'h%h !== 'hf", ir); end	// Vector No: 505
assert (op === 'hff) else begin fail = 1; $display("Error 2021: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2022: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2023: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// bfffffffffffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hbfffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 507
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2024: ir 'h%h !== 'hf", ir); end	// Vector No: 506
assert (op === 'hf8) else begin fail = 1; $display("Error 2025: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2026: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2027: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// bfffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hbfffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 508
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2028: ir 'h%h !== 'hf", ir); end	// Vector No: 507
assert (op === 'hf8) else begin fail = 1; $display("Error 2029: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2030: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2031: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 7fffffffffffffff:0:0:7:ff:0:fffff:
//------------------------

#2;
word <= 'h7fffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 509
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 2032: ir 'h%h !== 'h7", ir); end	// Vector No: 508
assert (op === 'hff) else begin fail = 1; $display("Error 2033: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2034: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2035: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 7fffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'h7fffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 510
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2036: ir 'h%h !== 'hf", ir); end	// Vector No: 509
assert (op === 'hff) else begin fail = 1; $display("Error 2037: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2038: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 2039: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 7fffffffffffffff:1:0:7:f8:0:07fff:
//------------------------

#2;
word <= 'h7fffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 511
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 2040: ir 'h%h !== 'h7", ir); end	// Vector No: 510
assert (op === 'hf8) else begin fail = 1; $display("Error 2041: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2042: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2043: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 7fffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'h7fffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 512
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 2044: ir 'h%h !== 'hf", ir); end	// Vector No: 511
assert (op === 'hf8) else begin fail = 1; $display("Error 2045: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2046: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 2047: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 0000000080000001:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 513
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2048: ir 'h%h !== 'h0", ir); end	// Vector No: 512
assert (op === 'h00) else begin fail = 1; $display("Error 2049: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2050: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2051: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000001:0:1:8:00:0:00001:
//------------------------

#2;
word <= 'h0000000080000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 514
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2052: ir 'h%h !== 'h8", ir); end	// Vector No: 513
assert (op === 'h00) else begin fail = 1; $display("Error 2053: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2054: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 2055: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000080000001:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 515
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2056: ir 'h%h !== 'h0", ir); end	// Vector No: 514
assert (op === 'h00) else begin fail = 1; $display("Error 2057: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2058: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2059: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000001:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 516
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2060: ir 'h%h !== 'h0", ir); end	// Vector No: 515
assert (op === 'h80) else begin fail = 1; $display("Error 2061: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2062: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2063: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000002:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000002;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 517
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2064: ir 'h%h !== 'h0", ir); end	// Vector No: 516
assert (op === 'h00) else begin fail = 1; $display("Error 2065: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2066: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2067: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000002:0:1:8:00:0:00002:
//------------------------

#2;
word <= 'h0000000080000002;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 518
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2068: ir 'h%h !== 'h8", ir); end	// Vector No: 517
assert (op === 'h00) else begin fail = 1; $display("Error 2069: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2070: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 2071: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000080000002:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000002;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 519
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2072: ir 'h%h !== 'h0", ir); end	// Vector No: 518
assert (op === 'h00) else begin fail = 1; $display("Error 2073: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2074: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2075: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000002:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000002;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 520
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2076: ir 'h%h !== 'h0", ir); end	// Vector No: 519
assert (op === 'h80) else begin fail = 1; $display("Error 2077: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2078: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2079: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000004:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000004;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 521
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2080: ir 'h%h !== 'h0", ir); end	// Vector No: 520
assert (op === 'h00) else begin fail = 1; $display("Error 2081: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2082: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2083: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000004:0:1:8:00:0:00004:
//------------------------

#2;
word <= 'h0000000080000004;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 522
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2084: ir 'h%h !== 'h8", ir); end	// Vector No: 521
assert (op === 'h00) else begin fail = 1; $display("Error 2085: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2086: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 2087: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000080000004:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000004;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 523
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2088: ir 'h%h !== 'h0", ir); end	// Vector No: 522
assert (op === 'h00) else begin fail = 1; $display("Error 2089: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2090: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2091: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000004:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000004;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 524
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2092: ir 'h%h !== 'h0", ir); end	// Vector No: 523
assert (op === 'h80) else begin fail = 1; $display("Error 2093: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2094: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2095: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000008:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000008;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 525
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2096: ir 'h%h !== 'h0", ir); end	// Vector No: 524
assert (op === 'h00) else begin fail = 1; $display("Error 2097: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2098: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2099: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000008:0:1:8:00:0:00008:
//------------------------

#2;
word <= 'h0000000080000008;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 526
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2100: ir 'h%h !== 'h8", ir); end	// Vector No: 525
assert (op === 'h00) else begin fail = 1; $display("Error 2101: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2102: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 2103: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000080000008:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000008;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 527
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2104: ir 'h%h !== 'h0", ir); end	// Vector No: 526
assert (op === 'h00) else begin fail = 1; $display("Error 2105: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2106: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2107: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000008:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000008;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 528
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2108: ir 'h%h !== 'h0", ir); end	// Vector No: 527
assert (op === 'h80) else begin fail = 1; $display("Error 2109: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2110: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2111: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000010:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 529
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2112: ir 'h%h !== 'h0", ir); end	// Vector No: 528
assert (op === 'h00) else begin fail = 1; $display("Error 2113: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2114: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2115: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000010:0:1:8:00:0:00010:
//------------------------

#2;
word <= 'h0000000080000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 530
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2116: ir 'h%h !== 'h8", ir); end	// Vector No: 529
assert (op === 'h00) else begin fail = 1; $display("Error 2117: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2118: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 2119: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000080000010:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 531
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2120: ir 'h%h !== 'h0", ir); end	// Vector No: 530
assert (op === 'h00) else begin fail = 1; $display("Error 2121: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2122: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2123: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000010:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 532
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2124: ir 'h%h !== 'h0", ir); end	// Vector No: 531
assert (op === 'h80) else begin fail = 1; $display("Error 2125: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2126: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2127: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000020:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000020;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 533
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2128: ir 'h%h !== 'h0", ir); end	// Vector No: 532
assert (op === 'h00) else begin fail = 1; $display("Error 2129: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2130: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2131: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000020:0:1:8:00:0:00020:
//------------------------

#2;
word <= 'h0000000080000020;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 534
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2132: ir 'h%h !== 'h8", ir); end	// Vector No: 533
assert (op === 'h00) else begin fail = 1; $display("Error 2133: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2134: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 2135: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000080000020:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000020;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 535
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2136: ir 'h%h !== 'h0", ir); end	// Vector No: 534
assert (op === 'h00) else begin fail = 1; $display("Error 2137: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2138: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2139: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000020:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000020;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 536
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2140: ir 'h%h !== 'h0", ir); end	// Vector No: 535
assert (op === 'h80) else begin fail = 1; $display("Error 2141: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2142: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2143: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000040:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000040;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 537
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2144: ir 'h%h !== 'h0", ir); end	// Vector No: 536
assert (op === 'h00) else begin fail = 1; $display("Error 2145: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2146: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2147: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000040:0:1:8:00:0:00040:
//------------------------

#2;
word <= 'h0000000080000040;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 538
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2148: ir 'h%h !== 'h8", ir); end	// Vector No: 537
assert (op === 'h00) else begin fail = 1; $display("Error 2149: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2150: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 2151: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000080000040:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000040;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 539
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2152: ir 'h%h !== 'h0", ir); end	// Vector No: 538
assert (op === 'h00) else begin fail = 1; $display("Error 2153: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2154: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2155: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000040:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000040;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 540
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2156: ir 'h%h !== 'h0", ir); end	// Vector No: 539
assert (op === 'h80) else begin fail = 1; $display("Error 2157: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2158: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2159: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000080:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000080;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 541
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2160: ir 'h%h !== 'h0", ir); end	// Vector No: 540
assert (op === 'h00) else begin fail = 1; $display("Error 2161: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2162: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2163: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000080:0:1:8:00:0:00080:
//------------------------

#2;
word <= 'h0000000080000080;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 542
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2164: ir 'h%h !== 'h8", ir); end	// Vector No: 541
assert (op === 'h00) else begin fail = 1; $display("Error 2165: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2166: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 2167: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000080000080:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000080;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 543
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2168: ir 'h%h !== 'h0", ir); end	// Vector No: 542
assert (op === 'h00) else begin fail = 1; $display("Error 2169: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2170: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2171: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000080:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000080;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 544
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2172: ir 'h%h !== 'h0", ir); end	// Vector No: 543
assert (op === 'h80) else begin fail = 1; $display("Error 2173: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2174: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2175: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000100:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 545
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2176: ir 'h%h !== 'h0", ir); end	// Vector No: 544
assert (op === 'h00) else begin fail = 1; $display("Error 2177: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2178: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2179: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000100:0:1:8:00:0:00100:
//------------------------

#2;
word <= 'h0000000080000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 546
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2180: ir 'h%h !== 'h8", ir); end	// Vector No: 545
assert (op === 'h00) else begin fail = 1; $display("Error 2181: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2182: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 2183: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000000080000100:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 547
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2184: ir 'h%h !== 'h0", ir); end	// Vector No: 546
assert (op === 'h00) else begin fail = 1; $display("Error 2185: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2186: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2187: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000100:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 548
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2188: ir 'h%h !== 'h0", ir); end	// Vector No: 547
assert (op === 'h80) else begin fail = 1; $display("Error 2189: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2190: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2191: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000200:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000200;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 549
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2192: ir 'h%h !== 'h0", ir); end	// Vector No: 548
assert (op === 'h00) else begin fail = 1; $display("Error 2193: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2194: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2195: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000200:0:1:8:00:0:00200:
//------------------------

#2;
word <= 'h0000000080000200;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 550
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2196: ir 'h%h !== 'h8", ir); end	// Vector No: 549
assert (op === 'h00) else begin fail = 1; $display("Error 2197: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2198: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 2199: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000000080000200:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000200;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 551
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2200: ir 'h%h !== 'h0", ir); end	// Vector No: 550
assert (op === 'h00) else begin fail = 1; $display("Error 2201: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2202: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2203: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000200:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000200;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 552
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2204: ir 'h%h !== 'h0", ir); end	// Vector No: 551
assert (op === 'h80) else begin fail = 1; $display("Error 2205: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2206: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2207: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000400:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000400;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 553
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2208: ir 'h%h !== 'h0", ir); end	// Vector No: 552
assert (op === 'h00) else begin fail = 1; $display("Error 2209: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2210: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2211: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000400:0:1:8:00:0:00400:
//------------------------

#2;
word <= 'h0000000080000400;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 554
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2212: ir 'h%h !== 'h8", ir); end	// Vector No: 553
assert (op === 'h00) else begin fail = 1; $display("Error 2213: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2214: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 2215: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000000080000400:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000400;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 555
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2216: ir 'h%h !== 'h0", ir); end	// Vector No: 554
assert (op === 'h00) else begin fail = 1; $display("Error 2217: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2218: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2219: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000400:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000400;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 556
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2220: ir 'h%h !== 'h0", ir); end	// Vector No: 555
assert (op === 'h80) else begin fail = 1; $display("Error 2221: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2222: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2223: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000800:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000800;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 557
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2224: ir 'h%h !== 'h0", ir); end	// Vector No: 556
assert (op === 'h00) else begin fail = 1; $display("Error 2225: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2226: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2227: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000800:0:1:8:00:0:00800:
//------------------------

#2;
word <= 'h0000000080000800;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 558
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2228: ir 'h%h !== 'h8", ir); end	// Vector No: 557
assert (op === 'h00) else begin fail = 1; $display("Error 2229: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2230: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 2231: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000000080000800:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080000800;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 559
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2232: ir 'h%h !== 'h0", ir); end	// Vector No: 558
assert (op === 'h00) else begin fail = 1; $display("Error 2233: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2234: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2235: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080000800:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000000080000800;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 560
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2236: ir 'h%h !== 'h0", ir); end	// Vector No: 559
assert (op === 'h80) else begin fail = 1; $display("Error 2237: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2238: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2239: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080001000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 561
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2240: ir 'h%h !== 'h0", ir); end	// Vector No: 560
assert (op === 'h00) else begin fail = 1; $display("Error 2241: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2242: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2243: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080001000:0:1:8:00:0:01000:
//------------------------

#2;
word <= 'h0000000080001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 562
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2244: ir 'h%h !== 'h8", ir); end	// Vector No: 561
assert (op === 'h00) else begin fail = 1; $display("Error 2245: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2246: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 2247: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000000080001000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 563
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2248: ir 'h%h !== 'h0", ir); end	// Vector No: 562
assert (op === 'h00) else begin fail = 1; $display("Error 2249: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2250: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2251: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080001000:1:1:0:80:0:00001:
//------------------------

#2;
word <= 'h0000000080001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 564
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2252: ir 'h%h !== 'h0", ir); end	// Vector No: 563
assert (op === 'h80) else begin fail = 1; $display("Error 2253: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2254: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 2255: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000080002000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080002000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 565
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2256: ir 'h%h !== 'h0", ir); end	// Vector No: 564
assert (op === 'h00) else begin fail = 1; $display("Error 2257: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2258: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2259: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080002000:0:1:8:00:0:02000:
//------------------------

#2;
word <= 'h0000000080002000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 566
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2260: ir 'h%h !== 'h8", ir); end	// Vector No: 565
assert (op === 'h00) else begin fail = 1; $display("Error 2261: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2262: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 2263: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000000080002000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080002000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 567
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2264: ir 'h%h !== 'h0", ir); end	// Vector No: 566
assert (op === 'h00) else begin fail = 1; $display("Error 2265: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2266: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2267: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080002000:1:1:0:80:0:00002:
//------------------------

#2;
word <= 'h0000000080002000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 568
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2268: ir 'h%h !== 'h0", ir); end	// Vector No: 567
assert (op === 'h80) else begin fail = 1; $display("Error 2269: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2270: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 2271: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000080004000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080004000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 569
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2272: ir 'h%h !== 'h0", ir); end	// Vector No: 568
assert (op === 'h00) else begin fail = 1; $display("Error 2273: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2274: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2275: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080004000:0:1:8:00:0:04000:
//------------------------

#2;
word <= 'h0000000080004000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 570
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2276: ir 'h%h !== 'h8", ir); end	// Vector No: 569
assert (op === 'h00) else begin fail = 1; $display("Error 2277: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2278: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 2279: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000000080004000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080004000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 571
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2280: ir 'h%h !== 'h0", ir); end	// Vector No: 570
assert (op === 'h00) else begin fail = 1; $display("Error 2281: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2282: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2283: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080004000:1:1:0:80:0:00004:
//------------------------

#2;
word <= 'h0000000080004000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 572
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2284: ir 'h%h !== 'h0", ir); end	// Vector No: 571
assert (op === 'h80) else begin fail = 1; $display("Error 2285: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2286: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 2287: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000080008000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080008000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 573
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2288: ir 'h%h !== 'h0", ir); end	// Vector No: 572
assert (op === 'h00) else begin fail = 1; $display("Error 2289: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2290: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2291: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080008000:0:1:8:00:0:08000:
//------------------------

#2;
word <= 'h0000000080008000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 574
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2292: ir 'h%h !== 'h8", ir); end	// Vector No: 573
assert (op === 'h00) else begin fail = 1; $display("Error 2293: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2294: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 2295: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000000080008000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080008000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 575
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2296: ir 'h%h !== 'h0", ir); end	// Vector No: 574
assert (op === 'h00) else begin fail = 1; $display("Error 2297: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2298: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2299: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080008000:1:1:0:80:0:00008:
//------------------------

#2;
word <= 'h0000000080008000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 576
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2300: ir 'h%h !== 'h0", ir); end	// Vector No: 575
assert (op === 'h80) else begin fail = 1; $display("Error 2301: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2302: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 2303: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000080010000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 577
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2304: ir 'h%h !== 'h0", ir); end	// Vector No: 576
assert (op === 'h00) else begin fail = 1; $display("Error 2305: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2306: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2307: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080010000:0:1:8:00:0:10000:
//------------------------

#2;
word <= 'h0000000080010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 578
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2308: ir 'h%h !== 'h8", ir); end	// Vector No: 577
assert (op === 'h00) else begin fail = 1; $display("Error 2309: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2310: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 2311: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0000000080010000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 579
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2312: ir 'h%h !== 'h0", ir); end	// Vector No: 578
assert (op === 'h00) else begin fail = 1; $display("Error 2313: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2314: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2315: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080010000:1:1:0:80:0:00010:
//------------------------

#2;
word <= 'h0000000080010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 580
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2316: ir 'h%h !== 'h0", ir); end	// Vector No: 579
assert (op === 'h80) else begin fail = 1; $display("Error 2317: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2318: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 2319: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000080020000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080020000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 581
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2320: ir 'h%h !== 'h0", ir); end	// Vector No: 580
assert (op === 'h00) else begin fail = 1; $display("Error 2321: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2322: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2323: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080020000:0:1:8:00:0:20000:
//------------------------

#2;
word <= 'h0000000080020000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 582
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2324: ir 'h%h !== 'h8", ir); end	// Vector No: 581
assert (op === 'h00) else begin fail = 1; $display("Error 2325: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2326: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 2327: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0000000080020000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080020000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 583
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2328: ir 'h%h !== 'h0", ir); end	// Vector No: 582
assert (op === 'h00) else begin fail = 1; $display("Error 2329: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2330: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2331: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080020000:1:1:0:80:0:00020:
//------------------------

#2;
word <= 'h0000000080020000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 584
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2332: ir 'h%h !== 'h0", ir); end	// Vector No: 583
assert (op === 'h80) else begin fail = 1; $display("Error 2333: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2334: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 2335: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000080040000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080040000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 585
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2336: ir 'h%h !== 'h0", ir); end	// Vector No: 584
assert (op === 'h00) else begin fail = 1; $display("Error 2337: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2338: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2339: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080040000:0:1:8:00:0:40000:
//------------------------

#2;
word <= 'h0000000080040000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 586
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2340: ir 'h%h !== 'h8", ir); end	// Vector No: 585
assert (op === 'h00) else begin fail = 1; $display("Error 2341: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2342: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 2343: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0000000080040000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080040000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 587
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2344: ir 'h%h !== 'h0", ir); end	// Vector No: 586
assert (op === 'h00) else begin fail = 1; $display("Error 2345: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2346: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2347: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080040000:1:1:0:80:0:00040:
//------------------------

#2;
word <= 'h0000000080040000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 588
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2348: ir 'h%h !== 'h0", ir); end	// Vector No: 587
assert (op === 'h80) else begin fail = 1; $display("Error 2349: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2350: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 2351: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000080080000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080080000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 589
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2352: ir 'h%h !== 'h0", ir); end	// Vector No: 588
assert (op === 'h00) else begin fail = 1; $display("Error 2353: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2354: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2355: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080080000:0:1:8:00:0:80000:
//------------------------

#2;
word <= 'h0000000080080000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 590
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2356: ir 'h%h !== 'h8", ir); end	// Vector No: 589
assert (op === 'h00) else begin fail = 1; $display("Error 2357: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2358: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 2359: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0000000080080000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080080000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 591
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2360: ir 'h%h !== 'h0", ir); end	// Vector No: 590
assert (op === 'h00) else begin fail = 1; $display("Error 2361: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2362: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2363: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080080000:1:1:0:80:0:00080:
//------------------------

#2;
word <= 'h0000000080080000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 592
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2364: ir 'h%h !== 'h0", ir); end	// Vector No: 591
assert (op === 'h80) else begin fail = 1; $display("Error 2365: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2366: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 2367: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000080100000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 593
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2368: ir 'h%h !== 'h0", ir); end	// Vector No: 592
assert (op === 'h00) else begin fail = 1; $display("Error 2369: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2370: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2371: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080100000:0:1:8:01:0:00000:
//------------------------

#2;
word <= 'h0000000080100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 594
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2372: ir 'h%h !== 'h8", ir); end	// Vector No: 593
assert (op === 'h01) else begin fail = 1; $display("Error 2373: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2374: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2375: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080100000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 595
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2376: ir 'h%h !== 'h0", ir); end	// Vector No: 594
assert (op === 'h00) else begin fail = 1; $display("Error 2377: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2378: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2379: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080100000:1:1:0:80:0:00100:
//------------------------

#2;
word <= 'h0000000080100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 596
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2380: ir 'h%h !== 'h0", ir); end	// Vector No: 595
assert (op === 'h80) else begin fail = 1; $display("Error 2381: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2382: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 2383: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000000080200000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080200000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 597
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2384: ir 'h%h !== 'h0", ir); end	// Vector No: 596
assert (op === 'h00) else begin fail = 1; $display("Error 2385: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2386: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2387: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080200000:0:1:8:02:0:00000:
//------------------------

#2;
word <= 'h0000000080200000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 598
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2388: ir 'h%h !== 'h8", ir); end	// Vector No: 597
assert (op === 'h02) else begin fail = 1; $display("Error 2389: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2390: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2391: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080200000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080200000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 599
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2392: ir 'h%h !== 'h0", ir); end	// Vector No: 598
assert (op === 'h00) else begin fail = 1; $display("Error 2393: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2394: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2395: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080200000:1:1:0:80:0:00200:
//------------------------

#2;
word <= 'h0000000080200000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 600
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2396: ir 'h%h !== 'h0", ir); end	// Vector No: 599
assert (op === 'h80) else begin fail = 1; $display("Error 2397: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2398: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 2399: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000000080400000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080400000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 601
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2400: ir 'h%h !== 'h0", ir); end	// Vector No: 600
assert (op === 'h00) else begin fail = 1; $display("Error 2401: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2402: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2403: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080400000:0:1:8:04:0:00000:
//------------------------

#2;
word <= 'h0000000080400000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 602
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2404: ir 'h%h !== 'h8", ir); end	// Vector No: 601
assert (op === 'h04) else begin fail = 1; $display("Error 2405: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2406: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2407: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080400000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080400000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 603
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2408: ir 'h%h !== 'h0", ir); end	// Vector No: 602
assert (op === 'h00) else begin fail = 1; $display("Error 2409: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2410: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2411: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080400000:1:1:0:80:0:00400:
//------------------------

#2;
word <= 'h0000000080400000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 604
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2412: ir 'h%h !== 'h0", ir); end	// Vector No: 603
assert (op === 'h80) else begin fail = 1; $display("Error 2413: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2414: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 2415: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000000080800000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080800000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 605
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2416: ir 'h%h !== 'h0", ir); end	// Vector No: 604
assert (op === 'h00) else begin fail = 1; $display("Error 2417: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2418: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2419: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080800000:0:1:8:08:0:00000:
//------------------------

#2;
word <= 'h0000000080800000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 606
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2420: ir 'h%h !== 'h8", ir); end	// Vector No: 605
assert (op === 'h08) else begin fail = 1; $display("Error 2421: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2422: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2423: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080800000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000080800000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 607
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2424: ir 'h%h !== 'h0", ir); end	// Vector No: 606
assert (op === 'h00) else begin fail = 1; $display("Error 2425: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2426: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2427: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000080800000:1:1:0:80:0:00800:
//------------------------

#2;
word <= 'h0000000080800000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 608
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2428: ir 'h%h !== 'h0", ir); end	// Vector No: 607
assert (op === 'h80) else begin fail = 1; $display("Error 2429: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2430: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 2431: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000000081000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000081000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 609
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2432: ir 'h%h !== 'h0", ir); end	// Vector No: 608
assert (op === 'h00) else begin fail = 1; $display("Error 2433: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2434: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2435: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000081000000:0:1:8:10:0:00000:
//------------------------

#2;
word <= 'h0000000081000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 610
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2436: ir 'h%h !== 'h8", ir); end	// Vector No: 609
assert (op === 'h10) else begin fail = 1; $display("Error 2437: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2438: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2439: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000081000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000081000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 611
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2440: ir 'h%h !== 'h0", ir); end	// Vector No: 610
assert (op === 'h00) else begin fail = 1; $display("Error 2441: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2442: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2443: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000081000000:1:1:0:80:0:01000:
//------------------------

#2;
word <= 'h0000000081000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 612
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2444: ir 'h%h !== 'h0", ir); end	// Vector No: 611
assert (op === 'h80) else begin fail = 1; $display("Error 2445: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2446: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 2447: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000000082000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000082000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 613
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2448: ir 'h%h !== 'h0", ir); end	// Vector No: 612
assert (op === 'h00) else begin fail = 1; $display("Error 2449: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2450: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2451: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000082000000:0:1:8:20:0:00000:
//------------------------

#2;
word <= 'h0000000082000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 614
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2452: ir 'h%h !== 'h8", ir); end	// Vector No: 613
assert (op === 'h20) else begin fail = 1; $display("Error 2453: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2454: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2455: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000082000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000082000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 615
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2456: ir 'h%h !== 'h0", ir); end	// Vector No: 614
assert (op === 'h00) else begin fail = 1; $display("Error 2457: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2458: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2459: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000082000000:1:1:0:80:0:02000:
//------------------------

#2;
word <= 'h0000000082000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 616
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2460: ir 'h%h !== 'h0", ir); end	// Vector No: 615
assert (op === 'h80) else begin fail = 1; $display("Error 2461: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2462: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 2463: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000000084000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000084000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 617
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2464: ir 'h%h !== 'h0", ir); end	// Vector No: 616
assert (op === 'h00) else begin fail = 1; $display("Error 2465: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2466: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2467: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000084000000:0:1:8:40:0:00000:
//------------------------

#2;
word <= 'h0000000084000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 618
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2468: ir 'h%h !== 'h8", ir); end	// Vector No: 617
assert (op === 'h40) else begin fail = 1; $display("Error 2469: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2470: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2471: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000084000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000084000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 619
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2472: ir 'h%h !== 'h0", ir); end	// Vector No: 618
assert (op === 'h00) else begin fail = 1; $display("Error 2473: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2474: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2475: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000084000000:1:1:0:80:0:04000:
//------------------------

#2;
word <= 'h0000000084000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 620
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2476: ir 'h%h !== 'h0", ir); end	// Vector No: 619
assert (op === 'h80) else begin fail = 1; $display("Error 2477: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2478: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 2479: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000000088000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000088000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 621
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2480: ir 'h%h !== 'h0", ir); end	// Vector No: 620
assert (op === 'h00) else begin fail = 1; $display("Error 2481: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2482: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2483: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000088000000:0:1:8:80:0:00000:
//------------------------

#2;
word <= 'h0000000088000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 622
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2484: ir 'h%h !== 'h8", ir); end	// Vector No: 621
assert (op === 'h80) else begin fail = 1; $display("Error 2485: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2486: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2487: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000088000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000088000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 623
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2488: ir 'h%h !== 'h0", ir); end	// Vector No: 622
assert (op === 'h00) else begin fail = 1; $display("Error 2489: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2490: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2491: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000088000000:1:1:0:88:0:00000:
//------------------------

#2;
word <= 'h0000000088000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 624
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2492: ir 'h%h !== 'h0", ir); end	// Vector No: 623
assert (op === 'h88) else begin fail = 1; $display("Error 2493: op 'h%h !== 'h88", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2494: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2495: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000090000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000090000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 625
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2496: ir 'h%h !== 'h0", ir); end	// Vector No: 624
assert (op === 'h00) else begin fail = 1; $display("Error 2497: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2498: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2499: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000090000000:0:1:9:00:0:00000:
//------------------------

#2;
word <= 'h0000000090000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 626
#2;

assert (ir === 'h9) else begin fail = 1; $display("Error 2500: ir 'h%h !== 'h9", ir); end	// Vector No: 625
assert (op === 'h00) else begin fail = 1; $display("Error 2501: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2502: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2503: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000090000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000090000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 627
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2504: ir 'h%h !== 'h0", ir); end	// Vector No: 626
assert (op === 'h00) else begin fail = 1; $display("Error 2505: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2506: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2507: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000090000000:1:1:0:90:0:00000:
//------------------------

#2;
word <= 'h0000000090000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 628
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2508: ir 'h%h !== 'h0", ir); end	// Vector No: 627
assert (op === 'h90) else begin fail = 1; $display("Error 2509: op 'h%h !== 'h90", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2510: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2511: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000a0000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h00000000a0000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 629
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2512: ir 'h%h !== 'h0", ir); end	// Vector No: 628
assert (op === 'h00) else begin fail = 1; $display("Error 2513: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2514: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2515: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000a0000000:0:1:a:00:0:00000:
//------------------------

#2;
word <= 'h00000000a0000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 630
#2;

assert (ir === 'ha) else begin fail = 1; $display("Error 2516: ir 'h%h !== 'ha", ir); end	// Vector No: 629
assert (op === 'h00) else begin fail = 1; $display("Error 2517: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2518: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2519: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000a0000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h00000000a0000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 631
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2520: ir 'h%h !== 'h0", ir); end	// Vector No: 630
assert (op === 'h00) else begin fail = 1; $display("Error 2521: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2522: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2523: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000a0000000:1:1:0:a0:0:00000:
//------------------------

#2;
word <= 'h00000000a0000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 632
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2524: ir 'h%h !== 'h0", ir); end	// Vector No: 631
assert (op === 'ha0) else begin fail = 1; $display("Error 2525: op 'h%h !== 'ha0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2526: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2527: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000c0000000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h00000000c0000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 633
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2528: ir 'h%h !== 'h0", ir); end	// Vector No: 632
assert (op === 'h00) else begin fail = 1; $display("Error 2529: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2530: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2531: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000c0000000:0:1:c:00:0:00000:
//------------------------

#2;
word <= 'h00000000c0000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 634
#2;

assert (ir === 'hc) else begin fail = 1; $display("Error 2532: ir 'h%h !== 'hc", ir); end	// Vector No: 633
assert (op === 'h00) else begin fail = 1; $display("Error 2533: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2534: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2535: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000c0000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h00000000c0000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 635
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2536: ir 'h%h !== 'h0", ir); end	// Vector No: 634
assert (op === 'h00) else begin fail = 1; $display("Error 2537: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2538: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2539: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00000000c0000000:1:1:0:c0:0:00000:
//------------------------

#2;
word <= 'h00000000c0000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 636
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2540: ir 'h%h !== 'h0", ir); end	// Vector No: 635
assert (op === 'hc0) else begin fail = 1; $display("Error 2541: op 'h%h !== 'hc0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2542: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2543: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000180000000:0:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000000180000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 637
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2544: ir 'h%h !== 'h0", ir); end	// Vector No: 636
assert (op === 'h00) else begin fail = 1; $display("Error 2545: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2546: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 2547: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000180000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000180000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 638
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2548: ir 'h%h !== 'h8", ir); end	// Vector No: 637
assert (op === 'h00) else begin fail = 1; $display("Error 2549: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2550: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2551: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000180000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000180000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 639
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2552: ir 'h%h !== 'h0", ir); end	// Vector No: 638
assert (op === 'h00) else begin fail = 1; $display("Error 2553: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2554: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2555: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000180000000:1:1:1:80:0:00000:
//------------------------

#2;
word <= 'h0000000180000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 640
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 2556: ir 'h%h !== 'h1", ir); end	// Vector No: 639
assert (op === 'h80) else begin fail = 1; $display("Error 2557: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2558: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2559: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000280000000:0:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000000280000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 641
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2560: ir 'h%h !== 'h0", ir); end	// Vector No: 640
assert (op === 'h00) else begin fail = 1; $display("Error 2561: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2562: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 2563: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000280000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000280000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 642
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2564: ir 'h%h !== 'h8", ir); end	// Vector No: 641
assert (op === 'h00) else begin fail = 1; $display("Error 2565: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2566: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2567: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000280000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000280000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 643
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2568: ir 'h%h !== 'h0", ir); end	// Vector No: 642
assert (op === 'h00) else begin fail = 1; $display("Error 2569: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2570: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2571: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000280000000:1:1:2:80:0:00000:
//------------------------

#2;
word <= 'h0000000280000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 644
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 2572: ir 'h%h !== 'h2", ir); end	// Vector No: 643
assert (op === 'h80) else begin fail = 1; $display("Error 2573: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2574: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2575: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000480000000:0:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000000480000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 645
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2576: ir 'h%h !== 'h0", ir); end	// Vector No: 644
assert (op === 'h00) else begin fail = 1; $display("Error 2577: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2578: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 2579: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000480000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000480000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 646
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2580: ir 'h%h !== 'h8", ir); end	// Vector No: 645
assert (op === 'h00) else begin fail = 1; $display("Error 2581: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2582: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2583: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000480000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000480000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 647
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2584: ir 'h%h !== 'h0", ir); end	// Vector No: 646
assert (op === 'h00) else begin fail = 1; $display("Error 2585: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2586: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2587: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000480000000:1:1:4:80:0:00000:
//------------------------

#2;
word <= 'h0000000480000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 648
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 2588: ir 'h%h !== 'h4", ir); end	// Vector No: 647
assert (op === 'h80) else begin fail = 1; $display("Error 2589: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2590: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2591: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000880000000:0:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000000880000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 649
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2592: ir 'h%h !== 'h0", ir); end	// Vector No: 648
assert (op === 'h00) else begin fail = 1; $display("Error 2593: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2594: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 2595: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000880000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000000880000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 650
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2596: ir 'h%h !== 'h8", ir); end	// Vector No: 649
assert (op === 'h00) else begin fail = 1; $display("Error 2597: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2598: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2599: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000880000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000880000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 651
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2600: ir 'h%h !== 'h0", ir); end	// Vector No: 650
assert (op === 'h00) else begin fail = 1; $display("Error 2601: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2602: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2603: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000880000000:1:1:8:80:0:00000:
//------------------------

#2;
word <= 'h0000000880000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 652
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2604: ir 'h%h !== 'h8", ir); end	// Vector No: 651
assert (op === 'h80) else begin fail = 1; $display("Error 2605: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2606: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2607: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001080000000:0:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000001080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 653
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2608: ir 'h%h !== 'h0", ir); end	// Vector No: 652
assert (op === 'h00) else begin fail = 1; $display("Error 2609: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2610: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 2611: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000001080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000001080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 654
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2612: ir 'h%h !== 'h8", ir); end	// Vector No: 653
assert (op === 'h00) else begin fail = 1; $display("Error 2613: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2614: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2615: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001080000000:1:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000001080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 655
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2616: ir 'h%h !== 'h0", ir); end	// Vector No: 654
assert (op === 'h00) else begin fail = 1; $display("Error 2617: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2618: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 2619: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000001080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000001080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 656
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2620: ir 'h%h !== 'h0", ir); end	// Vector No: 655
assert (op === 'h80) else begin fail = 1; $display("Error 2621: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2622: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2623: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002080000000:0:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000002080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 657
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2624: ir 'h%h !== 'h0", ir); end	// Vector No: 656
assert (op === 'h00) else begin fail = 1; $display("Error 2625: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2626: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 2627: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000002080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000002080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 658
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2628: ir 'h%h !== 'h8", ir); end	// Vector No: 657
assert (op === 'h00) else begin fail = 1; $display("Error 2629: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2630: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2631: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002080000000:1:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000002080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 659
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2632: ir 'h%h !== 'h0", ir); end	// Vector No: 658
assert (op === 'h00) else begin fail = 1; $display("Error 2633: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2634: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 2635: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000002080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000002080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 660
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2636: ir 'h%h !== 'h0", ir); end	// Vector No: 659
assert (op === 'h80) else begin fail = 1; $display("Error 2637: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2638: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2639: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004080000000:0:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000004080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 661
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2640: ir 'h%h !== 'h0", ir); end	// Vector No: 660
assert (op === 'h00) else begin fail = 1; $display("Error 2641: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2642: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 2643: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000004080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000004080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 662
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2644: ir 'h%h !== 'h8", ir); end	// Vector No: 661
assert (op === 'h00) else begin fail = 1; $display("Error 2645: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2646: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2647: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004080000000:1:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000004080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 663
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2648: ir 'h%h !== 'h0", ir); end	// Vector No: 662
assert (op === 'h00) else begin fail = 1; $display("Error 2649: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2650: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 2651: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000004080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000004080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 664
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2652: ir 'h%h !== 'h0", ir); end	// Vector No: 663
assert (op === 'h80) else begin fail = 1; $display("Error 2653: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2654: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2655: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008080000000:0:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000008080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 665
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2656: ir 'h%h !== 'h0", ir); end	// Vector No: 664
assert (op === 'h00) else begin fail = 1; $display("Error 2657: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2658: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 2659: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000008080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000008080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 666
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2660: ir 'h%h !== 'h8", ir); end	// Vector No: 665
assert (op === 'h00) else begin fail = 1; $display("Error 2661: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2662: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2663: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008080000000:1:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000008080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 667
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2664: ir 'h%h !== 'h0", ir); end	// Vector No: 666
assert (op === 'h00) else begin fail = 1; $display("Error 2665: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2666: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 2667: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000008080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000008080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 668
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2668: ir 'h%h !== 'h0", ir); end	// Vector No: 667
assert (op === 'h80) else begin fail = 1; $display("Error 2669: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2670: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2671: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010080000000:0:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000010080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 669
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2672: ir 'h%h !== 'h0", ir); end	// Vector No: 668
assert (op === 'h00) else begin fail = 1; $display("Error 2673: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2674: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 2675: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000010080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000010080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 670
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2676: ir 'h%h !== 'h8", ir); end	// Vector No: 669
assert (op === 'h00) else begin fail = 1; $display("Error 2677: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2678: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2679: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010080000000:1:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000010080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 671
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2680: ir 'h%h !== 'h0", ir); end	// Vector No: 670
assert (op === 'h00) else begin fail = 1; $display("Error 2681: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2682: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 2683: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000010080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000010080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 672
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2684: ir 'h%h !== 'h0", ir); end	// Vector No: 671
assert (op === 'h80) else begin fail = 1; $display("Error 2685: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2686: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2687: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020080000000:0:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000020080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 673
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2688: ir 'h%h !== 'h0", ir); end	// Vector No: 672
assert (op === 'h00) else begin fail = 1; $display("Error 2689: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2690: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 2691: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000020080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000020080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 674
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2692: ir 'h%h !== 'h8", ir); end	// Vector No: 673
assert (op === 'h00) else begin fail = 1; $display("Error 2693: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2694: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2695: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020080000000:1:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000020080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 675
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2696: ir 'h%h !== 'h0", ir); end	// Vector No: 674
assert (op === 'h00) else begin fail = 1; $display("Error 2697: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2698: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 2699: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000020080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000020080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 676
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2700: ir 'h%h !== 'h0", ir); end	// Vector No: 675
assert (op === 'h80) else begin fail = 1; $display("Error 2701: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2702: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2703: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040080000000:0:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000040080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 677
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2704: ir 'h%h !== 'h0", ir); end	// Vector No: 676
assert (op === 'h00) else begin fail = 1; $display("Error 2705: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2706: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 2707: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000040080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000040080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 678
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2708: ir 'h%h !== 'h8", ir); end	// Vector No: 677
assert (op === 'h00) else begin fail = 1; $display("Error 2709: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2710: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2711: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040080000000:1:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000040080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 679
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2712: ir 'h%h !== 'h0", ir); end	// Vector No: 678
assert (op === 'h00) else begin fail = 1; $display("Error 2713: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2714: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 2715: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000040080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000040080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 680
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2716: ir 'h%h !== 'h0", ir); end	// Vector No: 679
assert (op === 'h80) else begin fail = 1; $display("Error 2717: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2718: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2719: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080080000000:0:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000080080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 681
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2720: ir 'h%h !== 'h0", ir); end	// Vector No: 680
assert (op === 'h00) else begin fail = 1; $display("Error 2721: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2722: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 2723: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000080080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000080080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 682
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2724: ir 'h%h !== 'h8", ir); end	// Vector No: 681
assert (op === 'h00) else begin fail = 1; $display("Error 2725: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2726: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2727: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080080000000:1:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000080080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 683
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2728: ir 'h%h !== 'h0", ir); end	// Vector No: 682
assert (op === 'h00) else begin fail = 1; $display("Error 2729: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2730: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 2731: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000080080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000080080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 684
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2732: ir 'h%h !== 'h0", ir); end	// Vector No: 683
assert (op === 'h80) else begin fail = 1; $display("Error 2733: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2734: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2735: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100080000000:0:0:0:00:0:01000:
//------------------------

#2;
word <= 'h0000100080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 685
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2736: ir 'h%h !== 'h0", ir); end	// Vector No: 684
assert (op === 'h00) else begin fail = 1; $display("Error 2737: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2738: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 2739: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000100080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000100080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 686
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2740: ir 'h%h !== 'h8", ir); end	// Vector No: 685
assert (op === 'h00) else begin fail = 1; $display("Error 2741: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2742: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2743: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100080000000:1:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000100080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 687
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2744: ir 'h%h !== 'h0", ir); end	// Vector No: 686
assert (op === 'h00) else begin fail = 1; $display("Error 2745: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2746: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 2747: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000100080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000100080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 688
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2748: ir 'h%h !== 'h0", ir); end	// Vector No: 687
assert (op === 'h80) else begin fail = 1; $display("Error 2749: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2750: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2751: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200080000000:0:0:0:00:0:02000:
//------------------------

#2;
word <= 'h0000200080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 689
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2752: ir 'h%h !== 'h0", ir); end	// Vector No: 688
assert (op === 'h00) else begin fail = 1; $display("Error 2753: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2754: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 2755: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000200080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000200080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 690
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2756: ir 'h%h !== 'h8", ir); end	// Vector No: 689
assert (op === 'h00) else begin fail = 1; $display("Error 2757: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2758: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2759: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200080000000:1:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000200080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 691
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2760: ir 'h%h !== 'h0", ir); end	// Vector No: 690
assert (op === 'h00) else begin fail = 1; $display("Error 2761: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2762: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 2763: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000200080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000200080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 692
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2764: ir 'h%h !== 'h0", ir); end	// Vector No: 691
assert (op === 'h80) else begin fail = 1; $display("Error 2765: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2766: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2767: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400080000000:0:0:0:00:0:04000:
//------------------------

#2;
word <= 'h0000400080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 693
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2768: ir 'h%h !== 'h0", ir); end	// Vector No: 692
assert (op === 'h00) else begin fail = 1; $display("Error 2769: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2770: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 2771: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000400080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000400080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 694
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2772: ir 'h%h !== 'h8", ir); end	// Vector No: 693
assert (op === 'h00) else begin fail = 1; $display("Error 2773: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2774: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2775: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400080000000:1:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000400080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 695
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2776: ir 'h%h !== 'h0", ir); end	// Vector No: 694
assert (op === 'h00) else begin fail = 1; $display("Error 2777: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2778: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 2779: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000400080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000400080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 696
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2780: ir 'h%h !== 'h0", ir); end	// Vector No: 695
assert (op === 'h80) else begin fail = 1; $display("Error 2781: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2782: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2783: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800080000000:0:0:0:00:0:08000:
//------------------------

#2;
word <= 'h0000800080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 697
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2784: ir 'h%h !== 'h0", ir); end	// Vector No: 696
assert (op === 'h00) else begin fail = 1; $display("Error 2785: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2786: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 2787: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000800080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0000800080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 698
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2788: ir 'h%h !== 'h8", ir); end	// Vector No: 697
assert (op === 'h00) else begin fail = 1; $display("Error 2789: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2790: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2791: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800080000000:1:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000800080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 699
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2792: ir 'h%h !== 'h0", ir); end	// Vector No: 698
assert (op === 'h00) else begin fail = 1; $display("Error 2793: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2794: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 2795: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000800080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0000800080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 700
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2796: ir 'h%h !== 'h0", ir); end	// Vector No: 699
assert (op === 'h80) else begin fail = 1; $display("Error 2797: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2798: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2799: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000080000000:0:0:0:00:0:10000:
//------------------------

#2;
word <= 'h0001000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 701
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2800: ir 'h%h !== 'h0", ir); end	// Vector No: 700
assert (op === 'h00) else begin fail = 1; $display("Error 2801: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2802: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 2803: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0001000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0001000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 702
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2804: ir 'h%h !== 'h8", ir); end	// Vector No: 701
assert (op === 'h00) else begin fail = 1; $display("Error 2805: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2806: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2807: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000080000000:1:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0001000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 703
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2808: ir 'h%h !== 'h0", ir); end	// Vector No: 702
assert (op === 'h01) else begin fail = 1; $display("Error 2809: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2810: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2811: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0001000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 704
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2812: ir 'h%h !== 'h0", ir); end	// Vector No: 703
assert (op === 'h80) else begin fail = 1; $display("Error 2813: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2814: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2815: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000080000000:0:0:0:00:0:20000:
//------------------------

#2;
word <= 'h0002000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 705
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2816: ir 'h%h !== 'h0", ir); end	// Vector No: 704
assert (op === 'h00) else begin fail = 1; $display("Error 2817: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2818: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 2819: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0002000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0002000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 706
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2820: ir 'h%h !== 'h8", ir); end	// Vector No: 705
assert (op === 'h00) else begin fail = 1; $display("Error 2821: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2822: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2823: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000080000000:1:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0002000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 707
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2824: ir 'h%h !== 'h0", ir); end	// Vector No: 706
assert (op === 'h02) else begin fail = 1; $display("Error 2825: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2826: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2827: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0002000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 708
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2828: ir 'h%h !== 'h0", ir); end	// Vector No: 707
assert (op === 'h80) else begin fail = 1; $display("Error 2829: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2830: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2831: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000080000000:0:0:0:00:0:40000:
//------------------------

#2;
word <= 'h0004000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 709
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2832: ir 'h%h !== 'h0", ir); end	// Vector No: 708
assert (op === 'h00) else begin fail = 1; $display("Error 2833: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2834: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 2835: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0004000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0004000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 710
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2836: ir 'h%h !== 'h8", ir); end	// Vector No: 709
assert (op === 'h00) else begin fail = 1; $display("Error 2837: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2838: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2839: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000080000000:1:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0004000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 711
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2840: ir 'h%h !== 'h0", ir); end	// Vector No: 710
assert (op === 'h04) else begin fail = 1; $display("Error 2841: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2842: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2843: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0004000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 712
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2844: ir 'h%h !== 'h0", ir); end	// Vector No: 711
assert (op === 'h80) else begin fail = 1; $display("Error 2845: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2846: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2847: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000080000000:0:0:0:00:0:80000:
//------------------------

#2;
word <= 'h0008000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 713
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2848: ir 'h%h !== 'h0", ir); end	// Vector No: 712
assert (op === 'h00) else begin fail = 1; $display("Error 2849: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2850: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 2851: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0008000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0008000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 714
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2852: ir 'h%h !== 'h8", ir); end	// Vector No: 713
assert (op === 'h00) else begin fail = 1; $display("Error 2853: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2854: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2855: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000080000000:1:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0008000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 715
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2856: ir 'h%h !== 'h0", ir); end	// Vector No: 714
assert (op === 'h08) else begin fail = 1; $display("Error 2857: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2858: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2859: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0008000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 716
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2860: ir 'h%h !== 'h0", ir); end	// Vector No: 715
assert (op === 'h80) else begin fail = 1; $display("Error 2861: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2862: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2863: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000080000000:0:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0010000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 717
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2864: ir 'h%h !== 'h0", ir); end	// Vector No: 716
assert (op === 'h01) else begin fail = 1; $display("Error 2865: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2866: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2867: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0010000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 718
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2868: ir 'h%h !== 'h8", ir); end	// Vector No: 717
assert (op === 'h00) else begin fail = 1; $display("Error 2869: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2870: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2871: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000080000000:1:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0010000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 719
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2872: ir 'h%h !== 'h0", ir); end	// Vector No: 718
assert (op === 'h10) else begin fail = 1; $display("Error 2873: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2874: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2875: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0010000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 720
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2876: ir 'h%h !== 'h0", ir); end	// Vector No: 719
assert (op === 'h80) else begin fail = 1; $display("Error 2877: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2878: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2879: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000080000000:0:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0020000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 721
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2880: ir 'h%h !== 'h0", ir); end	// Vector No: 720
assert (op === 'h02) else begin fail = 1; $display("Error 2881: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2882: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2883: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0020000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 722
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2884: ir 'h%h !== 'h8", ir); end	// Vector No: 721
assert (op === 'h00) else begin fail = 1; $display("Error 2885: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2886: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2887: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000080000000:1:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0020000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 723
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2888: ir 'h%h !== 'h0", ir); end	// Vector No: 722
assert (op === 'h20) else begin fail = 1; $display("Error 2889: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2890: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2891: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0020000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 724
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2892: ir 'h%h !== 'h0", ir); end	// Vector No: 723
assert (op === 'h80) else begin fail = 1; $display("Error 2893: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2894: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2895: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000080000000:0:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0040000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 725
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2896: ir 'h%h !== 'h0", ir); end	// Vector No: 724
assert (op === 'h04) else begin fail = 1; $display("Error 2897: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2898: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2899: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0040000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 726
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2900: ir 'h%h !== 'h8", ir); end	// Vector No: 725
assert (op === 'h00) else begin fail = 1; $display("Error 2901: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2902: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2903: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000080000000:1:0:0:40:0:07000:
//------------------------

#2;
word <= 'h0040000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 727
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2904: ir 'h%h !== 'h0", ir); end	// Vector No: 726
assert (op === 'h40) else begin fail = 1; $display("Error 2905: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2906: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 2907: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0040000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0040000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 728
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2908: ir 'h%h !== 'h0", ir); end	// Vector No: 727
assert (op === 'h80) else begin fail = 1; $display("Error 2909: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2910: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2911: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000080000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 729
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2912: ir 'h%h !== 'h0", ir); end	// Vector No: 728
assert (op === 'h08) else begin fail = 1; $display("Error 2913: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2914: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2915: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0080000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 730
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2916: ir 'h%h !== 'h8", ir); end	// Vector No: 729
assert (op === 'h00) else begin fail = 1; $display("Error 2917: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2918: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2919: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000080000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 731
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2920: ir 'h%h !== 'h0", ir); end	// Vector No: 730
assert (op === 'h80) else begin fail = 1; $display("Error 2921: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2922: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2923: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 732
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2924: ir 'h%h !== 'h0", ir); end	// Vector No: 731
assert (op === 'h80) else begin fail = 1; $display("Error 2925: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2926: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2927: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000080000000:0:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0100000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 733
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2928: ir 'h%h !== 'h0", ir); end	// Vector No: 732
assert (op === 'h10) else begin fail = 1; $display("Error 2929: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2930: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2931: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0100000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 734
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2932: ir 'h%h !== 'h8", ir); end	// Vector No: 733
assert (op === 'h00) else begin fail = 1; $display("Error 2933: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2934: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2935: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000080000000:1:0:1:00:0:00000:
//------------------------

#2;
word <= 'h0100000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 735
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 2936: ir 'h%h !== 'h1", ir); end	// Vector No: 734
assert (op === 'h00) else begin fail = 1; $display("Error 2937: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2938: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2939: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0100000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 736
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2940: ir 'h%h !== 'h0", ir); end	// Vector No: 735
assert (op === 'h80) else begin fail = 1; $display("Error 2941: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2942: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2943: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000080000000:0:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0200000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 737
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2944: ir 'h%h !== 'h0", ir); end	// Vector No: 736
assert (op === 'h20) else begin fail = 1; $display("Error 2945: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2946: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2947: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0200000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 738
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2948: ir 'h%h !== 'h8", ir); end	// Vector No: 737
assert (op === 'h00) else begin fail = 1; $display("Error 2949: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2950: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2951: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000080000000:1:0:2:00:0:00000:
//------------------------

#2;
word <= 'h0200000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 739
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 2952: ir 'h%h !== 'h2", ir); end	// Vector No: 738
assert (op === 'h00) else begin fail = 1; $display("Error 2953: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2954: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2955: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0200000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 740
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2956: ir 'h%h !== 'h0", ir); end	// Vector No: 739
assert (op === 'h80) else begin fail = 1; $display("Error 2957: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2958: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2959: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000080000000:0:0:0:40:0:00000:
//------------------------

#2;
word <= 'h0400000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 741
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2960: ir 'h%h !== 'h0", ir); end	// Vector No: 740
assert (op === 'h40) else begin fail = 1; $display("Error 2961: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2962: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2963: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0400000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 742
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2964: ir 'h%h !== 'h8", ir); end	// Vector No: 741
assert (op === 'h00) else begin fail = 1; $display("Error 2965: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2966: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2967: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000080000000:1:0:4:00:0:00000:
//------------------------

#2;
word <= 'h0400000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 743
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 2968: ir 'h%h !== 'h4", ir); end	// Vector No: 742
assert (op === 'h00) else begin fail = 1; $display("Error 2969: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2970: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2971: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0400000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 744
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2972: ir 'h%h !== 'h0", ir); end	// Vector No: 743
assert (op === 'h80) else begin fail = 1; $display("Error 2973: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2974: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2975: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000080000000:0:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0800000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 745
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2976: ir 'h%h !== 'h0", ir); end	// Vector No: 744
assert (op === 'h80) else begin fail = 1; $display("Error 2977: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2978: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2979: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0800000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 746
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2980: ir 'h%h !== 'h8", ir); end	// Vector No: 745
assert (op === 'h00) else begin fail = 1; $display("Error 2981: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2982: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2983: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000080000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0800000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 747
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2984: ir 'h%h !== 'h0", ir); end	// Vector No: 746
assert (op === 'h00) else begin fail = 1; $display("Error 2985: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2986: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2987: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0800000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 748
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 2988: ir 'h%h !== 'h0", ir); end	// Vector No: 747
assert (op === 'h80) else begin fail = 1; $display("Error 2989: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2990: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2991: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000080000000:0:0:1:00:0:00000:
//------------------------

#2;
word <= 'h1000000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 749
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 2992: ir 'h%h !== 'h1", ir); end	// Vector No: 748
assert (op === 'h00) else begin fail = 1; $display("Error 2993: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2994: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2995: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h1000000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 750
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 2996: ir 'h%h !== 'h8", ir); end	// Vector No: 749
assert (op === 'h00) else begin fail = 1; $display("Error 2997: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 2998: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 2999: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000080000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h1000000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 751
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3000: ir 'h%h !== 'h0", ir); end	// Vector No: 750
assert (op === 'h00) else begin fail = 1; $display("Error 3001: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3002: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3003: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h1000000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 752
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3004: ir 'h%h !== 'h0", ir); end	// Vector No: 751
assert (op === 'h80) else begin fail = 1; $display("Error 3005: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3006: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3007: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000080000000:0:0:2:00:0:00000:
//------------------------

#2;
word <= 'h2000000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 753
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 3008: ir 'h%h !== 'h2", ir); end	// Vector No: 752
assert (op === 'h00) else begin fail = 1; $display("Error 3009: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3010: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3011: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h2000000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 754
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3012: ir 'h%h !== 'h8", ir); end	// Vector No: 753
assert (op === 'h00) else begin fail = 1; $display("Error 3013: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3014: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3015: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000080000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h2000000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 755
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3016: ir 'h%h !== 'h0", ir); end	// Vector No: 754
assert (op === 'h00) else begin fail = 1; $display("Error 3017: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3018: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3019: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h2000000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 756
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3020: ir 'h%h !== 'h0", ir); end	// Vector No: 755
assert (op === 'h80) else begin fail = 1; $display("Error 3021: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3022: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3023: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000080000000:0:0:4:00:0:00000:
//------------------------

#2;
word <= 'h4000000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 757
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 3024: ir 'h%h !== 'h4", ir); end	// Vector No: 756
assert (op === 'h00) else begin fail = 1; $display("Error 3025: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3026: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3027: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h4000000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 758
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3028: ir 'h%h !== 'h8", ir); end	// Vector No: 757
assert (op === 'h00) else begin fail = 1; $display("Error 3029: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3030: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3031: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000080000000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h4000000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 759
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3032: ir 'h%h !== 'h0", ir); end	// Vector No: 758
assert (op === 'h00) else begin fail = 1; $display("Error 3033: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3034: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3035: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h4000000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 760
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3036: ir 'h%h !== 'h0", ir); end	// Vector No: 759
assert (op === 'h80) else begin fail = 1; $display("Error 3037: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3038: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3039: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000080000000:0:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 761
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3040: ir 'h%h !== 'h8", ir); end	// Vector No: 760
assert (op === 'h00) else begin fail = 1; $display("Error 3041: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3042: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3043: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 762
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3044: ir 'h%h !== 'h8", ir); end	// Vector No: 761
assert (op === 'h00) else begin fail = 1; $display("Error 3045: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3046: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3047: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000080000000:1:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 763
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3048: ir 'h%h !== 'h8", ir); end	// Vector No: 762
assert (op === 'h00) else begin fail = 1; $display("Error 3049: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3050: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3051: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h8000000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 764
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3052: ir 'h%h !== 'h0", ir); end	// Vector No: 763
assert (op === 'h80) else begin fail = 1; $display("Error 3053: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3054: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3055: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000001:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 765
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3056: ir 'h%h !== 'h0", ir); end	// Vector No: 764
assert (op === 'h08) else begin fail = 1; $display("Error 3057: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3058: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3059: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000001:0:1:0:00:0:00001:
//------------------------

#2;
word <= 'h0080000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 766
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3060: ir 'h%h !== 'h0", ir); end	// Vector No: 765
assert (op === 'h00) else begin fail = 1; $display("Error 3061: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3062: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 3063: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0080000000000001:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 767
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3064: ir 'h%h !== 'h0", ir); end	// Vector No: 766
assert (op === 'h80) else begin fail = 1; $display("Error 3065: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3066: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3067: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000001:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 768
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3068: ir 'h%h !== 'h0", ir); end	// Vector No: 767
assert (op === 'h00) else begin fail = 1; $display("Error 3069: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3070: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3071: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000002:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000002;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 769
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3072: ir 'h%h !== 'h0", ir); end	// Vector No: 768
assert (op === 'h08) else begin fail = 1; $display("Error 3073: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3074: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3075: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000002:0:1:0:00:0:00002:
//------------------------

#2;
word <= 'h0080000000000002;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 770
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3076: ir 'h%h !== 'h0", ir); end	// Vector No: 769
assert (op === 'h00) else begin fail = 1; $display("Error 3077: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3078: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 3079: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0080000000000002:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000002;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 771
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3080: ir 'h%h !== 'h0", ir); end	// Vector No: 770
assert (op === 'h80) else begin fail = 1; $display("Error 3081: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3082: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3083: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000002:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000002;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 772
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3084: ir 'h%h !== 'h0", ir); end	// Vector No: 771
assert (op === 'h00) else begin fail = 1; $display("Error 3085: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3086: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3087: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000004:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000004;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 773
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3088: ir 'h%h !== 'h0", ir); end	// Vector No: 772
assert (op === 'h08) else begin fail = 1; $display("Error 3089: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3090: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3091: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000004:0:1:0:00:0:00004:
//------------------------

#2;
word <= 'h0080000000000004;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 774
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3092: ir 'h%h !== 'h0", ir); end	// Vector No: 773
assert (op === 'h00) else begin fail = 1; $display("Error 3093: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3094: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 3095: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0080000000000004:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000004;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 775
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3096: ir 'h%h !== 'h0", ir); end	// Vector No: 774
assert (op === 'h80) else begin fail = 1; $display("Error 3097: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3098: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3099: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000004:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000004;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 776
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3100: ir 'h%h !== 'h0", ir); end	// Vector No: 775
assert (op === 'h00) else begin fail = 1; $display("Error 3101: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3102: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3103: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000008:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000008;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 777
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3104: ir 'h%h !== 'h0", ir); end	// Vector No: 776
assert (op === 'h08) else begin fail = 1; $display("Error 3105: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3106: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3107: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000008:0:1:0:00:0:00008:
//------------------------

#2;
word <= 'h0080000000000008;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 778
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3108: ir 'h%h !== 'h0", ir); end	// Vector No: 777
assert (op === 'h00) else begin fail = 1; $display("Error 3109: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3110: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 3111: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0080000000000008:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000008;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 779
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3112: ir 'h%h !== 'h0", ir); end	// Vector No: 778
assert (op === 'h80) else begin fail = 1; $display("Error 3113: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3114: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3115: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000008:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000008;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 780
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3116: ir 'h%h !== 'h0", ir); end	// Vector No: 779
assert (op === 'h00) else begin fail = 1; $display("Error 3117: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3118: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3119: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000010:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 781
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3120: ir 'h%h !== 'h0", ir); end	// Vector No: 780
assert (op === 'h08) else begin fail = 1; $display("Error 3121: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3122: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3123: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000010:0:1:0:00:0:00010:
//------------------------

#2;
word <= 'h0080000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 782
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3124: ir 'h%h !== 'h0", ir); end	// Vector No: 781
assert (op === 'h00) else begin fail = 1; $display("Error 3125: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3126: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 3127: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0080000000000010:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 783
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3128: ir 'h%h !== 'h0", ir); end	// Vector No: 782
assert (op === 'h80) else begin fail = 1; $display("Error 3129: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3130: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3131: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000010:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 784
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3132: ir 'h%h !== 'h0", ir); end	// Vector No: 783
assert (op === 'h00) else begin fail = 1; $display("Error 3133: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3134: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3135: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000020:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000020;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 785
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3136: ir 'h%h !== 'h0", ir); end	// Vector No: 784
assert (op === 'h08) else begin fail = 1; $display("Error 3137: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3138: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3139: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000020:0:1:0:00:0:00020:
//------------------------

#2;
word <= 'h0080000000000020;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 786
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3140: ir 'h%h !== 'h0", ir); end	// Vector No: 785
assert (op === 'h00) else begin fail = 1; $display("Error 3141: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3142: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 3143: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0080000000000020:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000020;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 787
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3144: ir 'h%h !== 'h0", ir); end	// Vector No: 786
assert (op === 'h80) else begin fail = 1; $display("Error 3145: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3146: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3147: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000020:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000020;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 788
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3148: ir 'h%h !== 'h0", ir); end	// Vector No: 787
assert (op === 'h00) else begin fail = 1; $display("Error 3149: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3150: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3151: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000040:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000040;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 789
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3152: ir 'h%h !== 'h0", ir); end	// Vector No: 788
assert (op === 'h08) else begin fail = 1; $display("Error 3153: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3154: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3155: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000040:0:1:0:00:0:00040:
//------------------------

#2;
word <= 'h0080000000000040;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 790
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3156: ir 'h%h !== 'h0", ir); end	// Vector No: 789
assert (op === 'h00) else begin fail = 1; $display("Error 3157: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3158: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 3159: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0080000000000040:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000040;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 791
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3160: ir 'h%h !== 'h0", ir); end	// Vector No: 790
assert (op === 'h80) else begin fail = 1; $display("Error 3161: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3162: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3163: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000040:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000040;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 792
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3164: ir 'h%h !== 'h0", ir); end	// Vector No: 791
assert (op === 'h00) else begin fail = 1; $display("Error 3165: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3166: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3167: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000080:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000080;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 793
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3168: ir 'h%h !== 'h0", ir); end	// Vector No: 792
assert (op === 'h08) else begin fail = 1; $display("Error 3169: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3170: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3171: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000080:0:1:0:00:0:00080:
//------------------------

#2;
word <= 'h0080000000000080;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 794
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3172: ir 'h%h !== 'h0", ir); end	// Vector No: 793
assert (op === 'h00) else begin fail = 1; $display("Error 3173: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3174: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 3175: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0080000000000080:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000080;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 795
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3176: ir 'h%h !== 'h0", ir); end	// Vector No: 794
assert (op === 'h80) else begin fail = 1; $display("Error 3177: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3178: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3179: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000080:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000080;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 796
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3180: ir 'h%h !== 'h0", ir); end	// Vector No: 795
assert (op === 'h00) else begin fail = 1; $display("Error 3181: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3182: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3183: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000100:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 797
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3184: ir 'h%h !== 'h0", ir); end	// Vector No: 796
assert (op === 'h08) else begin fail = 1; $display("Error 3185: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3186: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3187: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000100:0:1:0:00:0:00100:
//------------------------

#2;
word <= 'h0080000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 798
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3188: ir 'h%h !== 'h0", ir); end	// Vector No: 797
assert (op === 'h00) else begin fail = 1; $display("Error 3189: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3190: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 3191: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0080000000000100:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 799
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3192: ir 'h%h !== 'h0", ir); end	// Vector No: 798
assert (op === 'h80) else begin fail = 1; $display("Error 3193: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3194: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3195: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000100:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 800
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3196: ir 'h%h !== 'h0", ir); end	// Vector No: 799
assert (op === 'h00) else begin fail = 1; $display("Error 3197: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3198: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3199: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000200:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000200;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 801
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3200: ir 'h%h !== 'h0", ir); end	// Vector No: 800
assert (op === 'h08) else begin fail = 1; $display("Error 3201: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3202: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3203: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000200:0:1:0:00:0:00200:
//------------------------

#2;
word <= 'h0080000000000200;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 802
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3204: ir 'h%h !== 'h0", ir); end	// Vector No: 801
assert (op === 'h00) else begin fail = 1; $display("Error 3205: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3206: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 3207: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0080000000000200:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000200;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 803
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3208: ir 'h%h !== 'h0", ir); end	// Vector No: 802
assert (op === 'h80) else begin fail = 1; $display("Error 3209: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3210: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3211: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000200:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000200;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 804
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3212: ir 'h%h !== 'h0", ir); end	// Vector No: 803
assert (op === 'h00) else begin fail = 1; $display("Error 3213: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3214: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3215: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000400:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000400;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 805
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3216: ir 'h%h !== 'h0", ir); end	// Vector No: 804
assert (op === 'h08) else begin fail = 1; $display("Error 3217: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3218: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3219: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000400:0:1:0:00:0:00400:
//------------------------

#2;
word <= 'h0080000000000400;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 806
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3220: ir 'h%h !== 'h0", ir); end	// Vector No: 805
assert (op === 'h00) else begin fail = 1; $display("Error 3221: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3222: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 3223: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0080000000000400:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000400;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 807
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3224: ir 'h%h !== 'h0", ir); end	// Vector No: 806
assert (op === 'h80) else begin fail = 1; $display("Error 3225: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3226: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3227: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000400:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000400;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 808
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3228: ir 'h%h !== 'h0", ir); end	// Vector No: 807
assert (op === 'h00) else begin fail = 1; $display("Error 3229: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3230: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3231: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000800:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000000800;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 809
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3232: ir 'h%h !== 'h0", ir); end	// Vector No: 808
assert (op === 'h08) else begin fail = 1; $display("Error 3233: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3234: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3235: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000800:0:1:0:00:0:00800:
//------------------------

#2;
word <= 'h0080000000000800;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 810
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3236: ir 'h%h !== 'h0", ir); end	// Vector No: 809
assert (op === 'h00) else begin fail = 1; $display("Error 3237: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3238: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 3239: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0080000000000800:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000000800;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 811
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3240: ir 'h%h !== 'h0", ir); end	// Vector No: 810
assert (op === 'h80) else begin fail = 1; $display("Error 3241: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3242: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3243: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000000800:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000000000800;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 812
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3244: ir 'h%h !== 'h0", ir); end	// Vector No: 811
assert (op === 'h00) else begin fail = 1; $display("Error 3245: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3246: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3247: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000001000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 813
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3248: ir 'h%h !== 'h0", ir); end	// Vector No: 812
assert (op === 'h08) else begin fail = 1; $display("Error 3249: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3250: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3251: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000001000:0:1:0:00:0:01000:
//------------------------

#2;
word <= 'h0080000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 814
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3252: ir 'h%h !== 'h0", ir); end	// Vector No: 813
assert (op === 'h00) else begin fail = 1; $display("Error 3253: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3254: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 3255: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0080000000001000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 815
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3256: ir 'h%h !== 'h0", ir); end	// Vector No: 814
assert (op === 'h80) else begin fail = 1; $display("Error 3257: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3258: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3259: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000001000:1:1:0:00:0:00001:
//------------------------

#2;
word <= 'h0080000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 816
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3260: ir 'h%h !== 'h0", ir); end	// Vector No: 815
assert (op === 'h00) else begin fail = 1; $display("Error 3261: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3262: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 3263: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0080000000002000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000002000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 817
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3264: ir 'h%h !== 'h0", ir); end	// Vector No: 816
assert (op === 'h08) else begin fail = 1; $display("Error 3265: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3266: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3267: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000002000:0:1:0:00:0:02000:
//------------------------

#2;
word <= 'h0080000000002000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 818
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3268: ir 'h%h !== 'h0", ir); end	// Vector No: 817
assert (op === 'h00) else begin fail = 1; $display("Error 3269: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3270: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 3271: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0080000000002000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000002000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 819
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3272: ir 'h%h !== 'h0", ir); end	// Vector No: 818
assert (op === 'h80) else begin fail = 1; $display("Error 3273: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3274: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3275: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000002000:1:1:0:00:0:00002:
//------------------------

#2;
word <= 'h0080000000002000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 820
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3276: ir 'h%h !== 'h0", ir); end	// Vector No: 819
assert (op === 'h00) else begin fail = 1; $display("Error 3277: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3278: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 3279: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0080000000004000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000004000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 821
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3280: ir 'h%h !== 'h0", ir); end	// Vector No: 820
assert (op === 'h08) else begin fail = 1; $display("Error 3281: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3282: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3283: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000004000:0:1:0:00:0:04000:
//------------------------

#2;
word <= 'h0080000000004000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 822
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3284: ir 'h%h !== 'h0", ir); end	// Vector No: 821
assert (op === 'h00) else begin fail = 1; $display("Error 3285: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3286: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 3287: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0080000000004000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000004000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 823
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3288: ir 'h%h !== 'h0", ir); end	// Vector No: 822
assert (op === 'h80) else begin fail = 1; $display("Error 3289: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3290: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3291: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000004000:1:1:0:00:0:00004:
//------------------------

#2;
word <= 'h0080000000004000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 824
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3292: ir 'h%h !== 'h0", ir); end	// Vector No: 823
assert (op === 'h00) else begin fail = 1; $display("Error 3293: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3294: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 3295: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0080000000008000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000008000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 825
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3296: ir 'h%h !== 'h0", ir); end	// Vector No: 824
assert (op === 'h08) else begin fail = 1; $display("Error 3297: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3298: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3299: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000008000:0:1:0:00:0:08000:
//------------------------

#2;
word <= 'h0080000000008000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 826
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3300: ir 'h%h !== 'h0", ir); end	// Vector No: 825
assert (op === 'h00) else begin fail = 1; $display("Error 3301: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3302: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 3303: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0080000000008000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000008000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 827
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3304: ir 'h%h !== 'h0", ir); end	// Vector No: 826
assert (op === 'h80) else begin fail = 1; $display("Error 3305: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3306: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3307: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000008000:1:1:0:00:0:00008:
//------------------------

#2;
word <= 'h0080000000008000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 828
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3308: ir 'h%h !== 'h0", ir); end	// Vector No: 827
assert (op === 'h00) else begin fail = 1; $display("Error 3309: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3310: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 3311: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0080000000010000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 829
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3312: ir 'h%h !== 'h0", ir); end	// Vector No: 828
assert (op === 'h08) else begin fail = 1; $display("Error 3313: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3314: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3315: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000010000:0:1:0:00:0:10000:
//------------------------

#2;
word <= 'h0080000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 830
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3316: ir 'h%h !== 'h0", ir); end	// Vector No: 829
assert (op === 'h00) else begin fail = 1; $display("Error 3317: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3318: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 3319: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0080000000010000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 831
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3320: ir 'h%h !== 'h0", ir); end	// Vector No: 830
assert (op === 'h80) else begin fail = 1; $display("Error 3321: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3322: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3323: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000010000:1:1:0:00:0:00010:
//------------------------

#2;
word <= 'h0080000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 832
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3324: ir 'h%h !== 'h0", ir); end	// Vector No: 831
assert (op === 'h00) else begin fail = 1; $display("Error 3325: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3326: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 3327: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0080000000020000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000020000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 833
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3328: ir 'h%h !== 'h0", ir); end	// Vector No: 832
assert (op === 'h08) else begin fail = 1; $display("Error 3329: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3330: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3331: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000020000:0:1:0:00:0:20000:
//------------------------

#2;
word <= 'h0080000000020000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 834
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3332: ir 'h%h !== 'h0", ir); end	// Vector No: 833
assert (op === 'h00) else begin fail = 1; $display("Error 3333: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3334: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 3335: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0080000000020000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000020000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 835
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3336: ir 'h%h !== 'h0", ir); end	// Vector No: 834
assert (op === 'h80) else begin fail = 1; $display("Error 3337: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3338: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3339: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000020000:1:1:0:00:0:00020:
//------------------------

#2;
word <= 'h0080000000020000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 836
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3340: ir 'h%h !== 'h0", ir); end	// Vector No: 835
assert (op === 'h00) else begin fail = 1; $display("Error 3341: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3342: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 3343: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0080000000040000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000040000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 837
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3344: ir 'h%h !== 'h0", ir); end	// Vector No: 836
assert (op === 'h08) else begin fail = 1; $display("Error 3345: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3346: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3347: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000040000:0:1:0:00:0:40000:
//------------------------

#2;
word <= 'h0080000000040000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 838
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3348: ir 'h%h !== 'h0", ir); end	// Vector No: 837
assert (op === 'h00) else begin fail = 1; $display("Error 3349: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3350: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 3351: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0080000000040000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000040000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 839
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3352: ir 'h%h !== 'h0", ir); end	// Vector No: 838
assert (op === 'h80) else begin fail = 1; $display("Error 3353: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3354: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3355: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000040000:1:1:0:00:0:00040:
//------------------------

#2;
word <= 'h0080000000040000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 840
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3356: ir 'h%h !== 'h0", ir); end	// Vector No: 839
assert (op === 'h00) else begin fail = 1; $display("Error 3357: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3358: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 3359: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0080000000080000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000080000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 841
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3360: ir 'h%h !== 'h0", ir); end	// Vector No: 840
assert (op === 'h08) else begin fail = 1; $display("Error 3361: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3362: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3363: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000080000:0:1:0:00:0:80000:
//------------------------

#2;
word <= 'h0080000000080000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 842
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3364: ir 'h%h !== 'h0", ir); end	// Vector No: 841
assert (op === 'h00) else begin fail = 1; $display("Error 3365: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3366: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 3367: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0080000000080000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000080000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 843
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3368: ir 'h%h !== 'h0", ir); end	// Vector No: 842
assert (op === 'h80) else begin fail = 1; $display("Error 3369: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3370: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3371: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000080000:1:1:0:00:0:00080:
//------------------------

#2;
word <= 'h0080000000080000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 844
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3372: ir 'h%h !== 'h0", ir); end	// Vector No: 843
assert (op === 'h00) else begin fail = 1; $display("Error 3373: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3374: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 3375: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0080000000100000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 845
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3376: ir 'h%h !== 'h0", ir); end	// Vector No: 844
assert (op === 'h08) else begin fail = 1; $display("Error 3377: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3378: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3379: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000100000:0:1:0:01:0:00000:
//------------------------

#2;
word <= 'h0080000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 846
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3380: ir 'h%h !== 'h0", ir); end	// Vector No: 845
assert (op === 'h01) else begin fail = 1; $display("Error 3381: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3382: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3383: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000100000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 847
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3384: ir 'h%h !== 'h0", ir); end	// Vector No: 846
assert (op === 'h80) else begin fail = 1; $display("Error 3385: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3386: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3387: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000100000:1:1:0:00:0:00100:
//------------------------

#2;
word <= 'h0080000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 848
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3388: ir 'h%h !== 'h0", ir); end	// Vector No: 847
assert (op === 'h00) else begin fail = 1; $display("Error 3389: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3390: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 3391: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0080000000200000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000200000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 849
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3392: ir 'h%h !== 'h0", ir); end	// Vector No: 848
assert (op === 'h08) else begin fail = 1; $display("Error 3393: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3394: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3395: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000200000:0:1:0:02:0:00000:
//------------------------

#2;
word <= 'h0080000000200000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 850
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3396: ir 'h%h !== 'h0", ir); end	// Vector No: 849
assert (op === 'h02) else begin fail = 1; $display("Error 3397: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3398: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3399: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000200000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000200000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 851
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3400: ir 'h%h !== 'h0", ir); end	// Vector No: 850
assert (op === 'h80) else begin fail = 1; $display("Error 3401: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3402: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3403: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000200000:1:1:0:00:0:00200:
//------------------------

#2;
word <= 'h0080000000200000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 852
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3404: ir 'h%h !== 'h0", ir); end	// Vector No: 851
assert (op === 'h00) else begin fail = 1; $display("Error 3405: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3406: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 3407: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0080000000400000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000400000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 853
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3408: ir 'h%h !== 'h0", ir); end	// Vector No: 852
assert (op === 'h08) else begin fail = 1; $display("Error 3409: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3410: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3411: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000400000:0:1:0:04:0:00000:
//------------------------

#2;
word <= 'h0080000000400000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 854
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3412: ir 'h%h !== 'h0", ir); end	// Vector No: 853
assert (op === 'h04) else begin fail = 1; $display("Error 3413: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3414: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3415: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000400000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000400000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 855
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3416: ir 'h%h !== 'h0", ir); end	// Vector No: 854
assert (op === 'h80) else begin fail = 1; $display("Error 3417: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3418: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3419: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000400000:1:1:0:00:0:00400:
//------------------------

#2;
word <= 'h0080000000400000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 856
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3420: ir 'h%h !== 'h0", ir); end	// Vector No: 855
assert (op === 'h00) else begin fail = 1; $display("Error 3421: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3422: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 3423: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0080000000800000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000800000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 857
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3424: ir 'h%h !== 'h0", ir); end	// Vector No: 856
assert (op === 'h08) else begin fail = 1; $display("Error 3425: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3426: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3427: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000800000:0:1:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000000800000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 858
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3428: ir 'h%h !== 'h0", ir); end	// Vector No: 857
assert (op === 'h08) else begin fail = 1; $display("Error 3429: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3430: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3431: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000800000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000000800000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 859
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3432: ir 'h%h !== 'h0", ir); end	// Vector No: 858
assert (op === 'h80) else begin fail = 1; $display("Error 3433: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3434: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3435: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000000800000:1:1:0:00:0:00800:
//------------------------

#2;
word <= 'h0080000000800000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 860
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3436: ir 'h%h !== 'h0", ir); end	// Vector No: 859
assert (op === 'h00) else begin fail = 1; $display("Error 3437: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3438: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 3439: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0080000001000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 861
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3440: ir 'h%h !== 'h0", ir); end	// Vector No: 860
assert (op === 'h08) else begin fail = 1; $display("Error 3441: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3442: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3443: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000001000000:0:1:0:10:0:00000:
//------------------------

#2;
word <= 'h0080000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 862
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3444: ir 'h%h !== 'h0", ir); end	// Vector No: 861
assert (op === 'h10) else begin fail = 1; $display("Error 3445: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3446: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3447: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000001000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 863
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3448: ir 'h%h !== 'h0", ir); end	// Vector No: 862
assert (op === 'h80) else begin fail = 1; $display("Error 3449: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3450: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3451: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000001000000:1:1:0:01:0:00000:
//------------------------

#2;
word <= 'h0080000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 864
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3452: ir 'h%h !== 'h0", ir); end	// Vector No: 863
assert (op === 'h01) else begin fail = 1; $display("Error 3453: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3454: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3455: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000002000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000002000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 865
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3456: ir 'h%h !== 'h0", ir); end	// Vector No: 864
assert (op === 'h08) else begin fail = 1; $display("Error 3457: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3458: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3459: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000002000000:0:1:0:20:0:00000:
//------------------------

#2;
word <= 'h0080000002000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 866
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3460: ir 'h%h !== 'h0", ir); end	// Vector No: 865
assert (op === 'h20) else begin fail = 1; $display("Error 3461: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3462: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3463: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000002000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000002000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 867
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3464: ir 'h%h !== 'h0", ir); end	// Vector No: 866
assert (op === 'h80) else begin fail = 1; $display("Error 3465: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3466: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3467: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000002000000:1:1:0:02:0:00000:
//------------------------

#2;
word <= 'h0080000002000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 868
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3468: ir 'h%h !== 'h0", ir); end	// Vector No: 867
assert (op === 'h02) else begin fail = 1; $display("Error 3469: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3470: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3471: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000004000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000004000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 869
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3472: ir 'h%h !== 'h0", ir); end	// Vector No: 868
assert (op === 'h08) else begin fail = 1; $display("Error 3473: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3474: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3475: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000004000000:0:1:0:40:0:00000:
//------------------------

#2;
word <= 'h0080000004000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 870
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3476: ir 'h%h !== 'h0", ir); end	// Vector No: 869
assert (op === 'h40) else begin fail = 1; $display("Error 3477: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3478: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3479: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000004000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000004000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 871
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3480: ir 'h%h !== 'h0", ir); end	// Vector No: 870
assert (op === 'h80) else begin fail = 1; $display("Error 3481: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3482: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3483: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000004000000:1:1:0:04:0:00000:
//------------------------

#2;
word <= 'h0080000004000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 872
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3484: ir 'h%h !== 'h0", ir); end	// Vector No: 871
assert (op === 'h04) else begin fail = 1; $display("Error 3485: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3486: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3487: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000008000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000008000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 873
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3488: ir 'h%h !== 'h0", ir); end	// Vector No: 872
assert (op === 'h08) else begin fail = 1; $display("Error 3489: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3490: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3491: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000008000000:0:1:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000008000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 874
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3492: ir 'h%h !== 'h0", ir); end	// Vector No: 873
assert (op === 'h80) else begin fail = 1; $display("Error 3493: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3494: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3495: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000008000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000008000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 875
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3496: ir 'h%h !== 'h0", ir); end	// Vector No: 874
assert (op === 'h80) else begin fail = 1; $display("Error 3497: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3498: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3499: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000008000000:1:1:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000008000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 876
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3500: ir 'h%h !== 'h0", ir); end	// Vector No: 875
assert (op === 'h08) else begin fail = 1; $display("Error 3501: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3502: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3503: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000010000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 877
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3504: ir 'h%h !== 'h0", ir); end	// Vector No: 876
assert (op === 'h08) else begin fail = 1; $display("Error 3505: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3506: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3507: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000010000000:0:1:1:00:0:00000:
//------------------------

#2;
word <= 'h0080000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 878
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 3508: ir 'h%h !== 'h1", ir); end	// Vector No: 877
assert (op === 'h00) else begin fail = 1; $display("Error 3509: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3510: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3511: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000010000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 879
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3512: ir 'h%h !== 'h0", ir); end	// Vector No: 878
assert (op === 'h80) else begin fail = 1; $display("Error 3513: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3514: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3515: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000010000000:1:1:0:10:0:00000:
//------------------------

#2;
word <= 'h0080000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 880
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3516: ir 'h%h !== 'h0", ir); end	// Vector No: 879
assert (op === 'h10) else begin fail = 1; $display("Error 3517: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3518: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3519: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000020000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000020000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 881
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3520: ir 'h%h !== 'h0", ir); end	// Vector No: 880
assert (op === 'h08) else begin fail = 1; $display("Error 3521: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3522: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3523: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000020000000:0:1:2:00:0:00000:
//------------------------

#2;
word <= 'h0080000020000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 882
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 3524: ir 'h%h !== 'h2", ir); end	// Vector No: 881
assert (op === 'h00) else begin fail = 1; $display("Error 3525: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3526: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3527: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000020000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000020000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 883
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3528: ir 'h%h !== 'h0", ir); end	// Vector No: 882
assert (op === 'h80) else begin fail = 1; $display("Error 3529: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3530: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3531: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000020000000:1:1:0:20:0:00000:
//------------------------

#2;
word <= 'h0080000020000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 884
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3532: ir 'h%h !== 'h0", ir); end	// Vector No: 883
assert (op === 'h20) else begin fail = 1; $display("Error 3533: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3534: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3535: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000040000000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000040000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 885
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3536: ir 'h%h !== 'h0", ir); end	// Vector No: 884
assert (op === 'h08) else begin fail = 1; $display("Error 3537: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3538: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3539: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000040000000:0:1:4:00:0:00000:
//------------------------

#2;
word <= 'h0080000040000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 886
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 3540: ir 'h%h !== 'h4", ir); end	// Vector No: 885
assert (op === 'h00) else begin fail = 1; $display("Error 3541: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3542: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3543: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000040000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000040000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 887
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3544: ir 'h%h !== 'h0", ir); end	// Vector No: 886
assert (op === 'h80) else begin fail = 1; $display("Error 3545: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3546: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3547: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000040000000:1:1:0:40:0:07000:
//------------------------

#2;
word <= 'h0080000040000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 888
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3548: ir 'h%h !== 'h0", ir); end	// Vector No: 887
assert (op === 'h40) else begin fail = 1; $display("Error 3549: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3550: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 3551: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0080000100000000:0:0:0:08:0:00001:
//------------------------

#2;
word <= 'h0080000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 889
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3552: ir 'h%h !== 'h0", ir); end	// Vector No: 888
assert (op === 'h08) else begin fail = 1; $display("Error 3553: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3554: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 3555: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0080000100000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 890
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3556: ir 'h%h !== 'h0", ir); end	// Vector No: 889
assert (op === 'h00) else begin fail = 1; $display("Error 3557: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3558: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3559: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000100000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 891
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3560: ir 'h%h !== 'h0", ir); end	// Vector No: 890
assert (op === 'h80) else begin fail = 1; $display("Error 3561: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3562: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3563: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000100000000:1:1:1:00:0:00000:
//------------------------

#2;
word <= 'h0080000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 892
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 3564: ir 'h%h !== 'h1", ir); end	// Vector No: 891
assert (op === 'h00) else begin fail = 1; $display("Error 3565: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3566: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3567: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000200000000:0:0:0:08:0:00002:
//------------------------

#2;
word <= 'h0080000200000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 893
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3568: ir 'h%h !== 'h0", ir); end	// Vector No: 892
assert (op === 'h08) else begin fail = 1; $display("Error 3569: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3570: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 3571: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0080000200000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000200000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 894
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3572: ir 'h%h !== 'h0", ir); end	// Vector No: 893
assert (op === 'h00) else begin fail = 1; $display("Error 3573: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3574: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3575: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000200000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000200000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 895
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3576: ir 'h%h !== 'h0", ir); end	// Vector No: 894
assert (op === 'h80) else begin fail = 1; $display("Error 3577: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3578: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3579: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000200000000:1:1:2:00:0:00000:
//------------------------

#2;
word <= 'h0080000200000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 896
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 3580: ir 'h%h !== 'h2", ir); end	// Vector No: 895
assert (op === 'h00) else begin fail = 1; $display("Error 3581: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3582: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3583: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000400000000:0:0:0:08:0:00004:
//------------------------

#2;
word <= 'h0080000400000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 897
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3584: ir 'h%h !== 'h0", ir); end	// Vector No: 896
assert (op === 'h08) else begin fail = 1; $display("Error 3585: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3586: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 3587: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0080000400000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000400000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 898
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3588: ir 'h%h !== 'h0", ir); end	// Vector No: 897
assert (op === 'h00) else begin fail = 1; $display("Error 3589: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3590: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3591: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000400000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000400000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 899
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3592: ir 'h%h !== 'h0", ir); end	// Vector No: 898
assert (op === 'h80) else begin fail = 1; $display("Error 3593: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3594: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3595: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000400000000:1:1:4:00:0:00000:
//------------------------

#2;
word <= 'h0080000400000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 900
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 3596: ir 'h%h !== 'h4", ir); end	// Vector No: 899
assert (op === 'h00) else begin fail = 1; $display("Error 3597: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3598: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3599: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000800000000:0:0:0:08:0:00008:
//------------------------

#2;
word <= 'h0080000800000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 901
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3600: ir 'h%h !== 'h0", ir); end	// Vector No: 900
assert (op === 'h08) else begin fail = 1; $display("Error 3601: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3602: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 3603: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0080000800000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080000800000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 902
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3604: ir 'h%h !== 'h0", ir); end	// Vector No: 901
assert (op === 'h00) else begin fail = 1; $display("Error 3605: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3606: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3607: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000800000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000800000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 903
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3608: ir 'h%h !== 'h0", ir); end	// Vector No: 902
assert (op === 'h80) else begin fail = 1; $display("Error 3609: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3610: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3611: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000800000000:1:1:8:00:0:00000:
//------------------------

#2;
word <= 'h0080000800000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 904
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 3612: ir 'h%h !== 'h8", ir); end	// Vector No: 903
assert (op === 'h00) else begin fail = 1; $display("Error 3613: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3614: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3615: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080001000000000:0:0:0:08:0:00010:
//------------------------

#2;
word <= 'h0080001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 905
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3616: ir 'h%h !== 'h0", ir); end	// Vector No: 904
assert (op === 'h08) else begin fail = 1; $display("Error 3617: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3618: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 3619: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0080001000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 906
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3620: ir 'h%h !== 'h0", ir); end	// Vector No: 905
assert (op === 'h00) else begin fail = 1; $display("Error 3621: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3622: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3623: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080001000000000:1:0:0:80:0:00001:
//------------------------

#2;
word <= 'h0080001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 907
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3624: ir 'h%h !== 'h0", ir); end	// Vector No: 906
assert (op === 'h80) else begin fail = 1; $display("Error 3625: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3626: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 3627: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0080001000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 908
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3628: ir 'h%h !== 'h0", ir); end	// Vector No: 907
assert (op === 'h00) else begin fail = 1; $display("Error 3629: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3630: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3631: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080002000000000:0:0:0:08:0:00020:
//------------------------

#2;
word <= 'h0080002000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 909
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3632: ir 'h%h !== 'h0", ir); end	// Vector No: 908
assert (op === 'h08) else begin fail = 1; $display("Error 3633: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3634: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 3635: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0080002000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080002000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 910
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3636: ir 'h%h !== 'h0", ir); end	// Vector No: 909
assert (op === 'h00) else begin fail = 1; $display("Error 3637: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3638: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3639: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080002000000000:1:0:0:80:0:00002:
//------------------------

#2;
word <= 'h0080002000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 911
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3640: ir 'h%h !== 'h0", ir); end	// Vector No: 910
assert (op === 'h80) else begin fail = 1; $display("Error 3641: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3642: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 3643: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0080002000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080002000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 912
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3644: ir 'h%h !== 'h0", ir); end	// Vector No: 911
assert (op === 'h00) else begin fail = 1; $display("Error 3645: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3646: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3647: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080004000000000:0:0:0:08:0:00040:
//------------------------

#2;
word <= 'h0080004000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 913
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3648: ir 'h%h !== 'h0", ir); end	// Vector No: 912
assert (op === 'h08) else begin fail = 1; $display("Error 3649: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3650: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 3651: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0080004000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080004000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 914
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3652: ir 'h%h !== 'h0", ir); end	// Vector No: 913
assert (op === 'h00) else begin fail = 1; $display("Error 3653: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3654: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3655: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080004000000000:1:0:0:80:0:00004:
//------------------------

#2;
word <= 'h0080004000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 915
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3656: ir 'h%h !== 'h0", ir); end	// Vector No: 914
assert (op === 'h80) else begin fail = 1; $display("Error 3657: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3658: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 3659: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0080004000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080004000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 916
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3660: ir 'h%h !== 'h0", ir); end	// Vector No: 915
assert (op === 'h00) else begin fail = 1; $display("Error 3661: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3662: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3663: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080008000000000:0:0:0:08:0:00080:
//------------------------

#2;
word <= 'h0080008000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 917
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3664: ir 'h%h !== 'h0", ir); end	// Vector No: 916
assert (op === 'h08) else begin fail = 1; $display("Error 3665: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3666: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 3667: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0080008000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080008000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 918
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3668: ir 'h%h !== 'h0", ir); end	// Vector No: 917
assert (op === 'h00) else begin fail = 1; $display("Error 3669: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3670: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3671: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080008000000000:1:0:0:80:0:00008:
//------------------------

#2;
word <= 'h0080008000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 919
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3672: ir 'h%h !== 'h0", ir); end	// Vector No: 918
assert (op === 'h80) else begin fail = 1; $display("Error 3673: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3674: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 3675: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0080008000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080008000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 920
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3676: ir 'h%h !== 'h0", ir); end	// Vector No: 919
assert (op === 'h00) else begin fail = 1; $display("Error 3677: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3678: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3679: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080010000000000:0:0:0:08:0:00100:
//------------------------

#2;
word <= 'h0080010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 921
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3680: ir 'h%h !== 'h0", ir); end	// Vector No: 920
assert (op === 'h08) else begin fail = 1; $display("Error 3681: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3682: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 3683: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0080010000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 922
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3684: ir 'h%h !== 'h0", ir); end	// Vector No: 921
assert (op === 'h00) else begin fail = 1; $display("Error 3685: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3686: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3687: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080010000000000:1:0:0:80:0:00010:
//------------------------

#2;
word <= 'h0080010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 923
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3688: ir 'h%h !== 'h0", ir); end	// Vector No: 922
assert (op === 'h80) else begin fail = 1; $display("Error 3689: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3690: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 3691: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0080010000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 924
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3692: ir 'h%h !== 'h0", ir); end	// Vector No: 923
assert (op === 'h00) else begin fail = 1; $display("Error 3693: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3694: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3695: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080020000000000:0:0:0:08:0:00200:
//------------------------

#2;
word <= 'h0080020000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 925
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3696: ir 'h%h !== 'h0", ir); end	// Vector No: 924
assert (op === 'h08) else begin fail = 1; $display("Error 3697: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3698: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 3699: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0080020000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080020000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 926
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3700: ir 'h%h !== 'h0", ir); end	// Vector No: 925
assert (op === 'h00) else begin fail = 1; $display("Error 3701: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3702: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3703: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080020000000000:1:0:0:80:0:00020:
//------------------------

#2;
word <= 'h0080020000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 927
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3704: ir 'h%h !== 'h0", ir); end	// Vector No: 926
assert (op === 'h80) else begin fail = 1; $display("Error 3705: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3706: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 3707: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0080020000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080020000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 928
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3708: ir 'h%h !== 'h0", ir); end	// Vector No: 927
assert (op === 'h00) else begin fail = 1; $display("Error 3709: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3710: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3711: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080040000000000:0:0:0:08:0:00400:
//------------------------

#2;
word <= 'h0080040000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 929
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3712: ir 'h%h !== 'h0", ir); end	// Vector No: 928
assert (op === 'h08) else begin fail = 1; $display("Error 3713: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3714: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 3715: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0080040000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080040000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 930
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3716: ir 'h%h !== 'h0", ir); end	// Vector No: 929
assert (op === 'h00) else begin fail = 1; $display("Error 3717: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3718: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3719: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080040000000000:1:0:0:80:0:00040:
//------------------------

#2;
word <= 'h0080040000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 931
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3720: ir 'h%h !== 'h0", ir); end	// Vector No: 930
assert (op === 'h80) else begin fail = 1; $display("Error 3721: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3722: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 3723: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0080040000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080040000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 932
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3724: ir 'h%h !== 'h0", ir); end	// Vector No: 931
assert (op === 'h00) else begin fail = 1; $display("Error 3725: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3726: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3727: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080080000000000:0:0:0:08:0:00800:
//------------------------

#2;
word <= 'h0080080000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 933
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3728: ir 'h%h !== 'h0", ir); end	// Vector No: 932
assert (op === 'h08) else begin fail = 1; $display("Error 3729: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3730: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 3731: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0080080000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080080000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 934
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3732: ir 'h%h !== 'h0", ir); end	// Vector No: 933
assert (op === 'h00) else begin fail = 1; $display("Error 3733: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3734: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3735: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080080000000000:1:0:0:80:0:00080:
//------------------------

#2;
word <= 'h0080080000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 935
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3736: ir 'h%h !== 'h0", ir); end	// Vector No: 934
assert (op === 'h80) else begin fail = 1; $display("Error 3737: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3738: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 3739: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0080080000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080080000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 936
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3740: ir 'h%h !== 'h0", ir); end	// Vector No: 935
assert (op === 'h00) else begin fail = 1; $display("Error 3741: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3742: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3743: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080100000000000:0:0:0:08:0:01000:
//------------------------

#2;
word <= 'h0080100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 937
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3744: ir 'h%h !== 'h0", ir); end	// Vector No: 936
assert (op === 'h08) else begin fail = 1; $display("Error 3745: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3746: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 3747: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0080100000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 938
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3748: ir 'h%h !== 'h0", ir); end	// Vector No: 937
assert (op === 'h00) else begin fail = 1; $display("Error 3749: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3750: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3751: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080100000000000:1:0:0:80:0:00100:
//------------------------

#2;
word <= 'h0080100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 939
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3752: ir 'h%h !== 'h0", ir); end	// Vector No: 938
assert (op === 'h80) else begin fail = 1; $display("Error 3753: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3754: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 3755: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0080100000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 940
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3756: ir 'h%h !== 'h0", ir); end	// Vector No: 939
assert (op === 'h00) else begin fail = 1; $display("Error 3757: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3758: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3759: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080200000000000:0:0:0:08:0:02000:
//------------------------

#2;
word <= 'h0080200000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 941
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3760: ir 'h%h !== 'h0", ir); end	// Vector No: 940
assert (op === 'h08) else begin fail = 1; $display("Error 3761: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3762: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 3763: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0080200000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080200000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 942
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3764: ir 'h%h !== 'h0", ir); end	// Vector No: 941
assert (op === 'h00) else begin fail = 1; $display("Error 3765: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3766: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3767: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080200000000000:1:0:0:80:0:00200:
//------------------------

#2;
word <= 'h0080200000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 943
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3768: ir 'h%h !== 'h0", ir); end	// Vector No: 942
assert (op === 'h80) else begin fail = 1; $display("Error 3769: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3770: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 3771: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0080200000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080200000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 944
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3772: ir 'h%h !== 'h0", ir); end	// Vector No: 943
assert (op === 'h00) else begin fail = 1; $display("Error 3773: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3774: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3775: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080400000000000:0:0:0:08:0:04000:
//------------------------

#2;
word <= 'h0080400000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 945
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3776: ir 'h%h !== 'h0", ir); end	// Vector No: 944
assert (op === 'h08) else begin fail = 1; $display("Error 3777: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3778: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 3779: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0080400000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080400000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 946
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3780: ir 'h%h !== 'h0", ir); end	// Vector No: 945
assert (op === 'h00) else begin fail = 1; $display("Error 3781: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3782: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3783: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080400000000000:1:0:0:80:0:00400:
//------------------------

#2;
word <= 'h0080400000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 947
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3784: ir 'h%h !== 'h0", ir); end	// Vector No: 946
assert (op === 'h80) else begin fail = 1; $display("Error 3785: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3786: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 3787: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0080400000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080400000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 948
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3788: ir 'h%h !== 'h0", ir); end	// Vector No: 947
assert (op === 'h00) else begin fail = 1; $display("Error 3789: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3790: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3791: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080800000000000:0:0:0:08:0:08000:
//------------------------

#2;
word <= 'h0080800000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 949
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3792: ir 'h%h !== 'h0", ir); end	// Vector No: 948
assert (op === 'h08) else begin fail = 1; $display("Error 3793: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3794: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 3795: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0080800000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080800000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 950
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3796: ir 'h%h !== 'h0", ir); end	// Vector No: 949
assert (op === 'h00) else begin fail = 1; $display("Error 3797: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3798: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3799: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080800000000000:1:0:0:80:0:00800:
//------------------------

#2;
word <= 'h0080800000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 951
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3800: ir 'h%h !== 'h0", ir); end	// Vector No: 950
assert (op === 'h80) else begin fail = 1; $display("Error 3801: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3802: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 3803: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0080800000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0080800000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 952
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3804: ir 'h%h !== 'h0", ir); end	// Vector No: 951
assert (op === 'h00) else begin fail = 1; $display("Error 3805: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3806: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3807: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0081000000000000:0:0:0:08:0:10000:
//------------------------

#2;
word <= 'h0081000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 953
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3808: ir 'h%h !== 'h0", ir); end	// Vector No: 952
assert (op === 'h08) else begin fail = 1; $display("Error 3809: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3810: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 3811: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0081000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0081000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 954
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3812: ir 'h%h !== 'h0", ir); end	// Vector No: 953
assert (op === 'h00) else begin fail = 1; $display("Error 3813: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3814: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3815: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0081000000000000:1:0:0:80:0:01000:
//------------------------

#2;
word <= 'h0081000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 955
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3816: ir 'h%h !== 'h0", ir); end	// Vector No: 954
assert (op === 'h80) else begin fail = 1; $display("Error 3817: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3818: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 3819: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0081000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0081000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 956
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3820: ir 'h%h !== 'h0", ir); end	// Vector No: 955
assert (op === 'h00) else begin fail = 1; $display("Error 3821: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3822: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3823: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0082000000000000:0:0:0:08:0:20000:
//------------------------

#2;
word <= 'h0082000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 957
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3824: ir 'h%h !== 'h0", ir); end	// Vector No: 956
assert (op === 'h08) else begin fail = 1; $display("Error 3825: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3826: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 3827: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0082000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0082000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 958
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3828: ir 'h%h !== 'h0", ir); end	// Vector No: 957
assert (op === 'h00) else begin fail = 1; $display("Error 3829: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3830: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3831: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0082000000000000:1:0:0:80:0:02000:
//------------------------

#2;
word <= 'h0082000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 959
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3832: ir 'h%h !== 'h0", ir); end	// Vector No: 958
assert (op === 'h80) else begin fail = 1; $display("Error 3833: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3834: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 3835: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0082000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0082000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 960
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3836: ir 'h%h !== 'h0", ir); end	// Vector No: 959
assert (op === 'h00) else begin fail = 1; $display("Error 3837: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3838: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3839: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0084000000000000:0:0:0:08:0:40000:
//------------------------

#2;
word <= 'h0084000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 961
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3840: ir 'h%h !== 'h0", ir); end	// Vector No: 960
assert (op === 'h08) else begin fail = 1; $display("Error 3841: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3842: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 3843: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0084000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0084000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 962
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3844: ir 'h%h !== 'h0", ir); end	// Vector No: 961
assert (op === 'h00) else begin fail = 1; $display("Error 3845: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3846: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3847: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0084000000000000:1:0:0:80:0:04000:
//------------------------

#2;
word <= 'h0084000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 963
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3848: ir 'h%h !== 'h0", ir); end	// Vector No: 962
assert (op === 'h80) else begin fail = 1; $display("Error 3849: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3850: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 3851: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0084000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0084000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 964
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3852: ir 'h%h !== 'h0", ir); end	// Vector No: 963
assert (op === 'h00) else begin fail = 1; $display("Error 3853: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3854: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3855: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0088000000000000:0:0:0:08:0:80000:
//------------------------

#2;
word <= 'h0088000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 965
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3856: ir 'h%h !== 'h0", ir); end	// Vector No: 964
assert (op === 'h08) else begin fail = 1; $display("Error 3857: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3858: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 3859: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0088000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0088000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 966
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3860: ir 'h%h !== 'h0", ir); end	// Vector No: 965
assert (op === 'h00) else begin fail = 1; $display("Error 3861: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3862: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3863: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0088000000000000:1:0:0:88:0:00000:
//------------------------

#2;
word <= 'h0088000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 967
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3864: ir 'h%h !== 'h0", ir); end	// Vector No: 966
assert (op === 'h88) else begin fail = 1; $display("Error 3865: op 'h%h !== 'h88", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3866: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3867: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0088000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0088000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 968
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3868: ir 'h%h !== 'h0", ir); end	// Vector No: 967
assert (op === 'h00) else begin fail = 1; $display("Error 3869: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3870: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3871: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0090000000000000:0:0:0:09:0:00000:
//------------------------

#2;
word <= 'h0090000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 969
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3872: ir 'h%h !== 'h0", ir); end	// Vector No: 968
assert (op === 'h09) else begin fail = 1; $display("Error 3873: op 'h%h !== 'h09", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3874: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3875: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0090000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0090000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 970
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3876: ir 'h%h !== 'h0", ir); end	// Vector No: 969
assert (op === 'h00) else begin fail = 1; $display("Error 3877: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3878: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3879: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0090000000000000:1:0:0:90:0:00000:
//------------------------

#2;
word <= 'h0090000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 971
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3880: ir 'h%h !== 'h0", ir); end	// Vector No: 970
assert (op === 'h90) else begin fail = 1; $display("Error 3881: op 'h%h !== 'h90", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3882: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3883: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0090000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0090000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 972
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3884: ir 'h%h !== 'h0", ir); end	// Vector No: 971
assert (op === 'h00) else begin fail = 1; $display("Error 3885: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3886: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3887: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00a0000000000000:0:0:0:0a:0:00000:
//------------------------

#2;
word <= 'h00a0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 973
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3888: ir 'h%h !== 'h0", ir); end	// Vector No: 972
assert (op === 'h0a) else begin fail = 1; $display("Error 3889: op 'h%h !== 'h0a", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3890: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3891: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00a0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h00a0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 974
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3892: ir 'h%h !== 'h0", ir); end	// Vector No: 973
assert (op === 'h00) else begin fail = 1; $display("Error 3893: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3894: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3895: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00a0000000000000:1:0:0:a0:0:00000:
//------------------------

#2;
word <= 'h00a0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 975
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3896: ir 'h%h !== 'h0", ir); end	// Vector No: 974
assert (op === 'ha0) else begin fail = 1; $display("Error 3897: op 'h%h !== 'ha0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3898: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3899: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00a0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h00a0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 976
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3900: ir 'h%h !== 'h0", ir); end	// Vector No: 975
assert (op === 'h00) else begin fail = 1; $display("Error 3901: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3902: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3903: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00c0000000000000:0:0:0:0c:0:00000:
//------------------------

#2;
word <= 'h00c0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 977
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3904: ir 'h%h !== 'h0", ir); end	// Vector No: 976
assert (op === 'h0c) else begin fail = 1; $display("Error 3905: op 'h%h !== 'h0c", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3906: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3907: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00c0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h00c0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 978
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3908: ir 'h%h !== 'h0", ir); end	// Vector No: 977
assert (op === 'h00) else begin fail = 1; $display("Error 3909: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3910: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3911: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00c0000000000000:1:0:0:c0:0:00000:
//------------------------

#2;
word <= 'h00c0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 979
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3912: ir 'h%h !== 'h0", ir); end	// Vector No: 978
assert (op === 'hc0) else begin fail = 1; $display("Error 3913: op 'h%h !== 'hc0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3914: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3915: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 00c0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h00c0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 980
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3916: ir 'h%h !== 'h0", ir); end	// Vector No: 979
assert (op === 'h00) else begin fail = 1; $display("Error 3917: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3918: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3919: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0180000000000000:0:0:0:18:0:00000:
//------------------------

#2;
word <= 'h0180000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 981
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3920: ir 'h%h !== 'h0", ir); end	// Vector No: 980
assert (op === 'h18) else begin fail = 1; $display("Error 3921: op 'h%h !== 'h18", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3922: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3923: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0180000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0180000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 982
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3924: ir 'h%h !== 'h0", ir); end	// Vector No: 981
assert (op === 'h00) else begin fail = 1; $display("Error 3925: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3926: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3927: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0180000000000000:1:0:1:80:0:00000:
//------------------------

#2;
word <= 'h0180000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 983
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 3928: ir 'h%h !== 'h1", ir); end	// Vector No: 982
assert (op === 'h80) else begin fail = 1; $display("Error 3929: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3930: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3931: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0180000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0180000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 984
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3932: ir 'h%h !== 'h0", ir); end	// Vector No: 983
assert (op === 'h00) else begin fail = 1; $display("Error 3933: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3934: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3935: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0280000000000000:0:0:0:28:0:00000:
//------------------------

#2;
word <= 'h0280000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 985
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3936: ir 'h%h !== 'h0", ir); end	// Vector No: 984
assert (op === 'h28) else begin fail = 1; $display("Error 3937: op 'h%h !== 'h28", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3938: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3939: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0280000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0280000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 986
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3940: ir 'h%h !== 'h0", ir); end	// Vector No: 985
assert (op === 'h00) else begin fail = 1; $display("Error 3941: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3942: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3943: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0280000000000000:1:0:2:80:0:00000:
//------------------------

#2;
word <= 'h0280000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 987
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 3944: ir 'h%h !== 'h2", ir); end	// Vector No: 986
assert (op === 'h80) else begin fail = 1; $display("Error 3945: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3946: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3947: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0280000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0280000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 988
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3948: ir 'h%h !== 'h0", ir); end	// Vector No: 987
assert (op === 'h00) else begin fail = 1; $display("Error 3949: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3950: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3951: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0480000000000000:0:0:0:48:0:00000:
//------------------------

#2;
word <= 'h0480000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 989
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3952: ir 'h%h !== 'h0", ir); end	// Vector No: 988
assert (op === 'h48) else begin fail = 1; $display("Error 3953: op 'h%h !== 'h48", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3954: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3955: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0480000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0480000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 990
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3956: ir 'h%h !== 'h0", ir); end	// Vector No: 989
assert (op === 'h00) else begin fail = 1; $display("Error 3957: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3958: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3959: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0480000000000000:1:0:4:80:0:00000:
//------------------------

#2;
word <= 'h0480000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 991
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 3960: ir 'h%h !== 'h4", ir); end	// Vector No: 990
assert (op === 'h80) else begin fail = 1; $display("Error 3961: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3962: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3963: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0480000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0480000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 992
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3964: ir 'h%h !== 'h0", ir); end	// Vector No: 991
assert (op === 'h00) else begin fail = 1; $display("Error 3965: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3966: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3967: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0880000000000000:0:0:0:88:0:00000:
//------------------------

#2;
word <= 'h0880000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 993
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3968: ir 'h%h !== 'h0", ir); end	// Vector No: 992
assert (op === 'h88) else begin fail = 1; $display("Error 3969: op 'h%h !== 'h88", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3970: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3971: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0880000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0880000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 994
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3972: ir 'h%h !== 'h0", ir); end	// Vector No: 993
assert (op === 'h00) else begin fail = 1; $display("Error 3973: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3974: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3975: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0880000000000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0880000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 995
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3976: ir 'h%h !== 'h0", ir); end	// Vector No: 994
assert (op === 'h80) else begin fail = 1; $display("Error 3977: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3978: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3979: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0880000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h0880000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 996
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3980: ir 'h%h !== 'h0", ir); end	// Vector No: 995
assert (op === 'h00) else begin fail = 1; $display("Error 3981: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3982: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3983: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1080000000000000:0:0:1:08:0:00000:
//------------------------

#2;
word <= 'h1080000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 997
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 3984: ir 'h%h !== 'h1", ir); end	// Vector No: 996
assert (op === 'h08) else begin fail = 1; $display("Error 3985: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3986: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3987: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1080000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h1080000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 998
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3988: ir 'h%h !== 'h0", ir); end	// Vector No: 997
assert (op === 'h00) else begin fail = 1; $display("Error 3989: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3990: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3991: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1080000000000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h1080000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 999
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3992: ir 'h%h !== 'h0", ir); end	// Vector No: 998
assert (op === 'h80) else begin fail = 1; $display("Error 3993: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3994: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3995: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1080000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h1080000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1000
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 3996: ir 'h%h !== 'h0", ir); end	// Vector No: 999
assert (op === 'h00) else begin fail = 1; $display("Error 3997: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 3998: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 3999: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2080000000000000:0:0:2:08:0:00000:
//------------------------

#2;
word <= 'h2080000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1001
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 4000: ir 'h%h !== 'h2", ir); end	// Vector No: 1000
assert (op === 'h08) else begin fail = 1; $display("Error 4001: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4002: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4003: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2080000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h2080000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1002
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4004: ir 'h%h !== 'h0", ir); end	// Vector No: 1001
assert (op === 'h00) else begin fail = 1; $display("Error 4005: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4006: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4007: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2080000000000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h2080000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1003
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4008: ir 'h%h !== 'h0", ir); end	// Vector No: 1002
assert (op === 'h80) else begin fail = 1; $display("Error 4009: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4010: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4011: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2080000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h2080000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1004
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4012: ir 'h%h !== 'h0", ir); end	// Vector No: 1003
assert (op === 'h00) else begin fail = 1; $display("Error 4013: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4014: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4015: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4080000000000000:0:0:4:08:0:00000:
//------------------------

#2;
word <= 'h4080000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1005
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 4016: ir 'h%h !== 'h4", ir); end	// Vector No: 1004
assert (op === 'h08) else begin fail = 1; $display("Error 4017: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4018: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4019: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4080000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h4080000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1006
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4020: ir 'h%h !== 'h0", ir); end	// Vector No: 1005
assert (op === 'h00) else begin fail = 1; $display("Error 4021: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4022: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4023: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4080000000000000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h4080000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1007
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4024: ir 'h%h !== 'h0", ir); end	// Vector No: 1006
assert (op === 'h80) else begin fail = 1; $display("Error 4025: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4026: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4027: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4080000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h4080000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1008
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4028: ir 'h%h !== 'h0", ir); end	// Vector No: 1007
assert (op === 'h00) else begin fail = 1; $display("Error 4029: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4030: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4031: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8080000000000000:0:0:8:08:0:00000:
//------------------------

#2;
word <= 'h8080000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1009
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 4032: ir 'h%h !== 'h8", ir); end	// Vector No: 1008
assert (op === 'h08) else begin fail = 1; $display("Error 4033: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4034: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4035: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8080000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h8080000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1010
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4036: ir 'h%h !== 'h0", ir); end	// Vector No: 1009
assert (op === 'h00) else begin fail = 1; $display("Error 4037: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4038: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4039: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8080000000000000:1:0:8:80:0:00000:
//------------------------

#2;
word <= 'h8080000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1011
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 4040: ir 'h%h !== 'h8", ir); end	// Vector No: 1010
assert (op === 'h80) else begin fail = 1; $display("Error 4041: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4042: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4043: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8080000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h8080000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1012
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4044: ir 'h%h !== 'h0", ir); end	// Vector No: 1011
assert (op === 'h00) else begin fail = 1; $display("Error 4045: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4046: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4047: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00001:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1013
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4048: ir 'h%h !== 'h0", ir); end	// Vector No: 1012
assert (op === 'h00) else begin fail = 1; $display("Error 4049: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4050: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4051: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00001:0:1:0:00:1:00001:
//------------------------

#2;
word <= 'h0000000003f00001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1014
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4052: ir 'h%h !== 'h0", ir); end	// Vector No: 1013
assert (op === 'h00) else begin fail = 1; $display("Error 4053: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4054: extop 'h%h !== 1", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 4055: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000003f00001:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1015
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4056: ir 'h%h !== 'h0", ir); end	// Vector No: 1014
assert (op === 'h00) else begin fail = 1; $display("Error 4057: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4058: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4059: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00001:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1016
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4060: ir 'h%h !== 'h0", ir); end	// Vector No: 1015
assert (op === 'h03) else begin fail = 1; $display("Error 4061: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4062: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4063: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000001:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1017
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4064: ir 'h%h !== 'h0", ir); end	// Vector No: 1016
assert (op === 'h00) else begin fail = 1; $display("Error 4065: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4066: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4067: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000001:0:1:0:00:0:00001:
//------------------------

#2;
word <= 'h03f0000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1018
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4068: ir 'h%h !== 'h0", ir); end	// Vector No: 1017
assert (op === 'h00) else begin fail = 1; $display("Error 4069: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4070: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 4071: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 03f0000000000001:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1019
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4072: ir 'h%h !== 'h3", ir); end	// Vector No: 1018
assert (op === 'hf0) else begin fail = 1; $display("Error 4073: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4074: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4075: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000001:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1020
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4076: ir 'h%h !== 'h0", ir); end	// Vector No: 1019
assert (op === 'h00) else begin fail = 1; $display("Error 4077: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4078: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4079: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00002:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00002;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1021
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4080: ir 'h%h !== 'h0", ir); end	// Vector No: 1020
assert (op === 'h00) else begin fail = 1; $display("Error 4081: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4082: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4083: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00002:0:1:0:00:1:00002:
//------------------------

#2;
word <= 'h0000000003f00002;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1022
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4084: ir 'h%h !== 'h0", ir); end	// Vector No: 1021
assert (op === 'h00) else begin fail = 1; $display("Error 4085: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4086: extop 'h%h !== 1", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 4087: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000003f00002:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00002;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1023
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4088: ir 'h%h !== 'h0", ir); end	// Vector No: 1022
assert (op === 'h00) else begin fail = 1; $display("Error 4089: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4090: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4091: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00002:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00002;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1024
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4092: ir 'h%h !== 'h0", ir); end	// Vector No: 1023
assert (op === 'h03) else begin fail = 1; $display("Error 4093: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4094: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4095: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000002:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000002;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1025
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4096: ir 'h%h !== 'h0", ir); end	// Vector No: 1024
assert (op === 'h00) else begin fail = 1; $display("Error 4097: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4098: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4099: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000002:0:1:0:00:0:00002:
//------------------------

#2;
word <= 'h03f0000000000002;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1026
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4100: ir 'h%h !== 'h0", ir); end	// Vector No: 1025
assert (op === 'h00) else begin fail = 1; $display("Error 4101: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4102: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 4103: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 03f0000000000002:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000002;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1027
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4104: ir 'h%h !== 'h3", ir); end	// Vector No: 1026
assert (op === 'hf0) else begin fail = 1; $display("Error 4105: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4106: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4107: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000002:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000002;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1028
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4108: ir 'h%h !== 'h0", ir); end	// Vector No: 1027
assert (op === 'h00) else begin fail = 1; $display("Error 4109: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4110: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4111: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00004:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00004;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1029
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4112: ir 'h%h !== 'h0", ir); end	// Vector No: 1028
assert (op === 'h00) else begin fail = 1; $display("Error 4113: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4114: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4115: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00004:0:1:0:00:1:00004:
//------------------------

#2;
word <= 'h0000000003f00004;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1030
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4116: ir 'h%h !== 'h0", ir); end	// Vector No: 1029
assert (op === 'h00) else begin fail = 1; $display("Error 4117: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4118: extop 'h%h !== 1", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 4119: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000003f00004:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00004;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1031
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4120: ir 'h%h !== 'h0", ir); end	// Vector No: 1030
assert (op === 'h00) else begin fail = 1; $display("Error 4121: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4122: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4123: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00004:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00004;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1032
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4124: ir 'h%h !== 'h0", ir); end	// Vector No: 1031
assert (op === 'h03) else begin fail = 1; $display("Error 4125: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4126: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4127: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000004:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000004;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1033
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4128: ir 'h%h !== 'h0", ir); end	// Vector No: 1032
assert (op === 'h00) else begin fail = 1; $display("Error 4129: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4130: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4131: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000004:0:1:0:00:0:00004:
//------------------------

#2;
word <= 'h03f0000000000004;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1034
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4132: ir 'h%h !== 'h0", ir); end	// Vector No: 1033
assert (op === 'h00) else begin fail = 1; $display("Error 4133: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4134: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 4135: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 03f0000000000004:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000004;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1035
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4136: ir 'h%h !== 'h3", ir); end	// Vector No: 1034
assert (op === 'hf0) else begin fail = 1; $display("Error 4137: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4138: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4139: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000004:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000004;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1036
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4140: ir 'h%h !== 'h0", ir); end	// Vector No: 1035
assert (op === 'h00) else begin fail = 1; $display("Error 4141: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4142: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4143: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00008:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00008;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1037
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4144: ir 'h%h !== 'h0", ir); end	// Vector No: 1036
assert (op === 'h00) else begin fail = 1; $display("Error 4145: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4146: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4147: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00008:0:1:0:00:1:00008:
//------------------------

#2;
word <= 'h0000000003f00008;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1038
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4148: ir 'h%h !== 'h0", ir); end	// Vector No: 1037
assert (op === 'h00) else begin fail = 1; $display("Error 4149: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4150: extop 'h%h !== 1", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 4151: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000003f00008:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00008;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1039
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4152: ir 'h%h !== 'h0", ir); end	// Vector No: 1038
assert (op === 'h00) else begin fail = 1; $display("Error 4153: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4154: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4155: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00008:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00008;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1040
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4156: ir 'h%h !== 'h0", ir); end	// Vector No: 1039
assert (op === 'h03) else begin fail = 1; $display("Error 4157: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4158: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4159: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000008:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000008;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1041
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4160: ir 'h%h !== 'h0", ir); end	// Vector No: 1040
assert (op === 'h00) else begin fail = 1; $display("Error 4161: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4162: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4163: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000008:0:1:0:00:0:00008:
//------------------------

#2;
word <= 'h03f0000000000008;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1042
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4164: ir 'h%h !== 'h0", ir); end	// Vector No: 1041
assert (op === 'h00) else begin fail = 1; $display("Error 4165: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4166: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 4167: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 03f0000000000008:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000008;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1043
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4168: ir 'h%h !== 'h3", ir); end	// Vector No: 1042
assert (op === 'hf0) else begin fail = 1; $display("Error 4169: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4170: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4171: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000008:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000008;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1044
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4172: ir 'h%h !== 'h0", ir); end	// Vector No: 1043
assert (op === 'h00) else begin fail = 1; $display("Error 4173: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4174: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4175: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00010:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1045
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4176: ir 'h%h !== 'h0", ir); end	// Vector No: 1044
assert (op === 'h00) else begin fail = 1; $display("Error 4177: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4178: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4179: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00010:0:1:0:00:1:00010:
//------------------------

#2;
word <= 'h0000000003f00010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1046
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4180: ir 'h%h !== 'h0", ir); end	// Vector No: 1045
assert (op === 'h00) else begin fail = 1; $display("Error 4181: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4182: extop 'h%h !== 1", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 4183: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000003f00010:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1047
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4184: ir 'h%h !== 'h0", ir); end	// Vector No: 1046
assert (op === 'h00) else begin fail = 1; $display("Error 4185: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4186: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4187: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00010:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1048
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4188: ir 'h%h !== 'h0", ir); end	// Vector No: 1047
assert (op === 'h03) else begin fail = 1; $display("Error 4189: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4190: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4191: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000010:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1049
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4192: ir 'h%h !== 'h0", ir); end	// Vector No: 1048
assert (op === 'h00) else begin fail = 1; $display("Error 4193: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4194: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4195: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000010:0:1:0:00:0:00010:
//------------------------

#2;
word <= 'h03f0000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1050
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4196: ir 'h%h !== 'h0", ir); end	// Vector No: 1049
assert (op === 'h00) else begin fail = 1; $display("Error 4197: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4198: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 4199: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 03f0000000000010:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1051
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4200: ir 'h%h !== 'h3", ir); end	// Vector No: 1050
assert (op === 'hf0) else begin fail = 1; $display("Error 4201: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4202: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4203: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000010:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1052
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4204: ir 'h%h !== 'h0", ir); end	// Vector No: 1051
assert (op === 'h00) else begin fail = 1; $display("Error 4205: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4206: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4207: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00020:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00020;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1053
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4208: ir 'h%h !== 'h0", ir); end	// Vector No: 1052
assert (op === 'h00) else begin fail = 1; $display("Error 4209: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4210: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4211: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00020:0:1:0:00:1:00020:
//------------------------

#2;
word <= 'h0000000003f00020;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1054
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4212: ir 'h%h !== 'h0", ir); end	// Vector No: 1053
assert (op === 'h00) else begin fail = 1; $display("Error 4213: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4214: extop 'h%h !== 1", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 4215: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000003f00020:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00020;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1055
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4216: ir 'h%h !== 'h0", ir); end	// Vector No: 1054
assert (op === 'h00) else begin fail = 1; $display("Error 4217: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4218: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4219: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00020:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00020;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1056
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4220: ir 'h%h !== 'h0", ir); end	// Vector No: 1055
assert (op === 'h03) else begin fail = 1; $display("Error 4221: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4222: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4223: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000020:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000020;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1057
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4224: ir 'h%h !== 'h0", ir); end	// Vector No: 1056
assert (op === 'h00) else begin fail = 1; $display("Error 4225: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4226: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4227: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000020:0:1:0:00:0:00020:
//------------------------

#2;
word <= 'h03f0000000000020;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1058
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4228: ir 'h%h !== 'h0", ir); end	// Vector No: 1057
assert (op === 'h00) else begin fail = 1; $display("Error 4229: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4230: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 4231: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 03f0000000000020:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000020;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1059
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4232: ir 'h%h !== 'h3", ir); end	// Vector No: 1058
assert (op === 'hf0) else begin fail = 1; $display("Error 4233: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4234: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4235: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000020:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000020;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1060
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4236: ir 'h%h !== 'h0", ir); end	// Vector No: 1059
assert (op === 'h00) else begin fail = 1; $display("Error 4237: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4238: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4239: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00040:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00040;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1061
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4240: ir 'h%h !== 'h0", ir); end	// Vector No: 1060
assert (op === 'h00) else begin fail = 1; $display("Error 4241: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4242: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4243: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00040:0:1:0:00:1:00040:
//------------------------

#2;
word <= 'h0000000003f00040;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1062
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4244: ir 'h%h !== 'h0", ir); end	// Vector No: 1061
assert (op === 'h00) else begin fail = 1; $display("Error 4245: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4246: extop 'h%h !== 1", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 4247: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000003f00040:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00040;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1063
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4248: ir 'h%h !== 'h0", ir); end	// Vector No: 1062
assert (op === 'h00) else begin fail = 1; $display("Error 4249: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4250: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4251: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00040:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00040;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1064
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4252: ir 'h%h !== 'h0", ir); end	// Vector No: 1063
assert (op === 'h03) else begin fail = 1; $display("Error 4253: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4254: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4255: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000040:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000040;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1065
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4256: ir 'h%h !== 'h0", ir); end	// Vector No: 1064
assert (op === 'h00) else begin fail = 1; $display("Error 4257: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4258: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4259: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000040:0:1:0:00:0:00040:
//------------------------

#2;
word <= 'h03f0000000000040;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1066
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4260: ir 'h%h !== 'h0", ir); end	// Vector No: 1065
assert (op === 'h00) else begin fail = 1; $display("Error 4261: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4262: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 4263: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 03f0000000000040:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000040;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1067
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4264: ir 'h%h !== 'h3", ir); end	// Vector No: 1066
assert (op === 'hf0) else begin fail = 1; $display("Error 4265: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4266: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4267: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000040:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000040;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1068
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4268: ir 'h%h !== 'h0", ir); end	// Vector No: 1067
assert (op === 'h00) else begin fail = 1; $display("Error 4269: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4270: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4271: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00080:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00080;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1069
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4272: ir 'h%h !== 'h0", ir); end	// Vector No: 1068
assert (op === 'h00) else begin fail = 1; $display("Error 4273: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4274: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4275: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00080:0:1:0:00:1:00080:
//------------------------

#2;
word <= 'h0000000003f00080;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1070
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4276: ir 'h%h !== 'h0", ir); end	// Vector No: 1069
assert (op === 'h00) else begin fail = 1; $display("Error 4277: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4278: extop 'h%h !== 1", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 4279: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000003f00080:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00080;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1071
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4280: ir 'h%h !== 'h0", ir); end	// Vector No: 1070
assert (op === 'h00) else begin fail = 1; $display("Error 4281: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4282: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4283: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00080:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00080;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1072
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4284: ir 'h%h !== 'h0", ir); end	// Vector No: 1071
assert (op === 'h03) else begin fail = 1; $display("Error 4285: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4286: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4287: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000080:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000080;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1073
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4288: ir 'h%h !== 'h0", ir); end	// Vector No: 1072
assert (op === 'h00) else begin fail = 1; $display("Error 4289: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4290: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4291: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000080:0:1:0:00:0:00080:
//------------------------

#2;
word <= 'h03f0000000000080;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1074
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4292: ir 'h%h !== 'h0", ir); end	// Vector No: 1073
assert (op === 'h00) else begin fail = 1; $display("Error 4293: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4294: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 4295: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 03f0000000000080:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000080;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1075
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4296: ir 'h%h !== 'h3", ir); end	// Vector No: 1074
assert (op === 'hf0) else begin fail = 1; $display("Error 4297: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4298: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4299: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000080:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000080;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1076
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4300: ir 'h%h !== 'h0", ir); end	// Vector No: 1075
assert (op === 'h00) else begin fail = 1; $display("Error 4301: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4302: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4303: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00100:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1077
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4304: ir 'h%h !== 'h0", ir); end	// Vector No: 1076
assert (op === 'h00) else begin fail = 1; $display("Error 4305: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4306: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4307: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00100:0:1:0:00:1:00100:
//------------------------

#2;
word <= 'h0000000003f00100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1078
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4308: ir 'h%h !== 'h0", ir); end	// Vector No: 1077
assert (op === 'h00) else begin fail = 1; $display("Error 4309: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4310: extop 'h%h !== 1", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 4311: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000000003f00100:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1079
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4312: ir 'h%h !== 'h0", ir); end	// Vector No: 1078
assert (op === 'h00) else begin fail = 1; $display("Error 4313: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4314: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4315: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00100:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1080
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4316: ir 'h%h !== 'h0", ir); end	// Vector No: 1079
assert (op === 'h03) else begin fail = 1; $display("Error 4317: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4318: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4319: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000100:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1081
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4320: ir 'h%h !== 'h0", ir); end	// Vector No: 1080
assert (op === 'h00) else begin fail = 1; $display("Error 4321: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4322: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4323: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000100:0:1:0:00:0:00100:
//------------------------

#2;
word <= 'h03f0000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1082
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4324: ir 'h%h !== 'h0", ir); end	// Vector No: 1081
assert (op === 'h00) else begin fail = 1; $display("Error 4325: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4326: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 4327: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 03f0000000000100:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1083
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4328: ir 'h%h !== 'h3", ir); end	// Vector No: 1082
assert (op === 'hf0) else begin fail = 1; $display("Error 4329: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4330: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4331: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000100:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1084
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4332: ir 'h%h !== 'h0", ir); end	// Vector No: 1083
assert (op === 'h00) else begin fail = 1; $display("Error 4333: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4334: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4335: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00200:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00200;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1085
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4336: ir 'h%h !== 'h0", ir); end	// Vector No: 1084
assert (op === 'h00) else begin fail = 1; $display("Error 4337: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4338: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4339: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00200:0:1:0:00:1:00200:
//------------------------

#2;
word <= 'h0000000003f00200;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1086
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4340: ir 'h%h !== 'h0", ir); end	// Vector No: 1085
assert (op === 'h00) else begin fail = 1; $display("Error 4341: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4342: extop 'h%h !== 1", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 4343: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000000003f00200:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00200;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1087
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4344: ir 'h%h !== 'h0", ir); end	// Vector No: 1086
assert (op === 'h00) else begin fail = 1; $display("Error 4345: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4346: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4347: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00200:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00200;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1088
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4348: ir 'h%h !== 'h0", ir); end	// Vector No: 1087
assert (op === 'h03) else begin fail = 1; $display("Error 4349: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4350: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4351: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000200:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000200;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1089
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4352: ir 'h%h !== 'h0", ir); end	// Vector No: 1088
assert (op === 'h00) else begin fail = 1; $display("Error 4353: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4354: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4355: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000200:0:1:0:00:0:00200:
//------------------------

#2;
word <= 'h03f0000000000200;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1090
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4356: ir 'h%h !== 'h0", ir); end	// Vector No: 1089
assert (op === 'h00) else begin fail = 1; $display("Error 4357: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4358: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 4359: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 03f0000000000200:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000200;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1091
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4360: ir 'h%h !== 'h3", ir); end	// Vector No: 1090
assert (op === 'hf0) else begin fail = 1; $display("Error 4361: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4362: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4363: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000200:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000200;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1092
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4364: ir 'h%h !== 'h0", ir); end	// Vector No: 1091
assert (op === 'h00) else begin fail = 1; $display("Error 4365: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4366: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4367: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00400:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00400;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1093
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4368: ir 'h%h !== 'h0", ir); end	// Vector No: 1092
assert (op === 'h00) else begin fail = 1; $display("Error 4369: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4370: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4371: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00400:0:1:0:00:1:00400:
//------------------------

#2;
word <= 'h0000000003f00400;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1094
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4372: ir 'h%h !== 'h0", ir); end	// Vector No: 1093
assert (op === 'h00) else begin fail = 1; $display("Error 4373: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4374: extop 'h%h !== 1", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 4375: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000000003f00400:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00400;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1095
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4376: ir 'h%h !== 'h0", ir); end	// Vector No: 1094
assert (op === 'h00) else begin fail = 1; $display("Error 4377: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4378: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4379: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00400:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00400;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1096
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4380: ir 'h%h !== 'h0", ir); end	// Vector No: 1095
assert (op === 'h03) else begin fail = 1; $display("Error 4381: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4382: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4383: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000400:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000400;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1097
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4384: ir 'h%h !== 'h0", ir); end	// Vector No: 1096
assert (op === 'h00) else begin fail = 1; $display("Error 4385: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4386: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4387: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000400:0:1:0:00:0:00400:
//------------------------

#2;
word <= 'h03f0000000000400;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1098
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4388: ir 'h%h !== 'h0", ir); end	// Vector No: 1097
assert (op === 'h00) else begin fail = 1; $display("Error 4389: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4390: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 4391: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 03f0000000000400:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000400;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1099
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4392: ir 'h%h !== 'h3", ir); end	// Vector No: 1098
assert (op === 'hf0) else begin fail = 1; $display("Error 4393: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4394: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4395: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000400:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000400;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1100
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4396: ir 'h%h !== 'h0", ir); end	// Vector No: 1099
assert (op === 'h00) else begin fail = 1; $display("Error 4397: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4398: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4399: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00800:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00800;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1101
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4400: ir 'h%h !== 'h0", ir); end	// Vector No: 1100
assert (op === 'h00) else begin fail = 1; $display("Error 4401: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4402: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4403: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00800:0:1:0:00:1:00800:
//------------------------

#2;
word <= 'h0000000003f00800;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1102
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4404: ir 'h%h !== 'h0", ir); end	// Vector No: 1101
assert (op === 'h00) else begin fail = 1; $display("Error 4405: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4406: extop 'h%h !== 1", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 4407: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000000003f00800:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00800;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1103
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4408: ir 'h%h !== 'h0", ir); end	// Vector No: 1102
assert (op === 'h00) else begin fail = 1; $display("Error 4409: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4410: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4411: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00800:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00800;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1104
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4412: ir 'h%h !== 'h0", ir); end	// Vector No: 1103
assert (op === 'h03) else begin fail = 1; $display("Error 4413: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4414: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4415: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000800:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000800;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1105
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4416: ir 'h%h !== 'h0", ir); end	// Vector No: 1104
assert (op === 'h00) else begin fail = 1; $display("Error 4417: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4418: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4419: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000800:0:1:0:00:0:00800:
//------------------------

#2;
word <= 'h03f0000000000800;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1106
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4420: ir 'h%h !== 'h0", ir); end	// Vector No: 1105
assert (op === 'h00) else begin fail = 1; $display("Error 4421: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4422: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 4423: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 03f0000000000800:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000800;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1107
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4424: ir 'h%h !== 'h3", ir); end	// Vector No: 1106
assert (op === 'hf0) else begin fail = 1; $display("Error 4425: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4426: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4427: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000800:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000800;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1108
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4428: ir 'h%h !== 'h0", ir); end	// Vector No: 1107
assert (op === 'h00) else begin fail = 1; $display("Error 4429: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4430: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4431: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f01000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f01000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1109
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4432: ir 'h%h !== 'h0", ir); end	// Vector No: 1108
assert (op === 'h00) else begin fail = 1; $display("Error 4433: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4434: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4435: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f01000:0:1:0:01:1:01000:
//------------------------

#2;
word <= 'h0000000003f01000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1110
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4436: ir 'h%h !== 'h0", ir); end	// Vector No: 1109
assert (op === 'h01) else begin fail = 1; $display("Error 4437: op 'h%h !== 'h01", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4438: extop 'h%h !== 1", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 4439: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000000003f01000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f01000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1111
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4440: ir 'h%h !== 'h0", ir); end	// Vector No: 1110
assert (op === 'h00) else begin fail = 1; $display("Error 4441: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4442: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4443: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f01000:1:1:0:03:0:00f01:
//------------------------

#2;
word <= 'h0000000003f01000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1112
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4444: ir 'h%h !== 'h0", ir); end	// Vector No: 1111
assert (op === 'h03) else begin fail = 1; $display("Error 4445: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4446: extop 'h%h !== 0", extop); end
assert (addr === 'h00f01) else begin fail = 1; $display("Error 4447: addr 'h%h !== 'h00f01", addr); end
#2;
clk <= 0;

// 03f0000000001000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1113
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4448: ir 'h%h !== 'h0", ir); end	// Vector No: 1112
assert (op === 'h00) else begin fail = 1; $display("Error 4449: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4450: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4451: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000001000:0:1:0:00:0:01000:
//------------------------

#2;
word <= 'h03f0000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1114
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4452: ir 'h%h !== 'h0", ir); end	// Vector No: 1113
assert (op === 'h00) else begin fail = 1; $display("Error 4453: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4454: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 4455: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 03f0000000001000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1115
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4456: ir 'h%h !== 'h3", ir); end	// Vector No: 1114
assert (op === 'hf0) else begin fail = 1; $display("Error 4457: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4458: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4459: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000001000:1:1:0:00:0:00001:
//------------------------

#2;
word <= 'h03f0000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1116
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4460: ir 'h%h !== 'h0", ir); end	// Vector No: 1115
assert (op === 'h00) else begin fail = 1; $display("Error 4461: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4462: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 4463: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000003f02000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f02000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1117
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4464: ir 'h%h !== 'h0", ir); end	// Vector No: 1116
assert (op === 'h00) else begin fail = 1; $display("Error 4465: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4466: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4467: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f02000:0:1:0:02:1:02000:
//------------------------

#2;
word <= 'h0000000003f02000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1118
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4468: ir 'h%h !== 'h0", ir); end	// Vector No: 1117
assert (op === 'h02) else begin fail = 1; $display("Error 4469: op 'h%h !== 'h02", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4470: extop 'h%h !== 1", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 4471: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000000003f02000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f02000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1119
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4472: ir 'h%h !== 'h0", ir); end	// Vector No: 1118
assert (op === 'h00) else begin fail = 1; $display("Error 4473: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4474: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4475: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f02000:1:1:0:03:0:00f02:
//------------------------

#2;
word <= 'h0000000003f02000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1120
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4476: ir 'h%h !== 'h0", ir); end	// Vector No: 1119
assert (op === 'h03) else begin fail = 1; $display("Error 4477: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4478: extop 'h%h !== 0", extop); end
assert (addr === 'h00f02) else begin fail = 1; $display("Error 4479: addr 'h%h !== 'h00f02", addr); end
#2;
clk <= 0;

// 03f0000000002000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000002000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1121
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4480: ir 'h%h !== 'h0", ir); end	// Vector No: 1120
assert (op === 'h00) else begin fail = 1; $display("Error 4481: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4482: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4483: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000002000:0:1:0:00:0:02000:
//------------------------

#2;
word <= 'h03f0000000002000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1122
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4484: ir 'h%h !== 'h0", ir); end	// Vector No: 1121
assert (op === 'h00) else begin fail = 1; $display("Error 4485: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4486: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 4487: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 03f0000000002000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000002000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1123
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4488: ir 'h%h !== 'h3", ir); end	// Vector No: 1122
assert (op === 'hf0) else begin fail = 1; $display("Error 4489: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4490: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4491: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000002000:1:1:0:00:0:00002:
//------------------------

#2;
word <= 'h03f0000000002000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1124
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4492: ir 'h%h !== 'h0", ir); end	// Vector No: 1123
assert (op === 'h00) else begin fail = 1; $display("Error 4493: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4494: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 4495: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000003f04000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f04000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1125
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4496: ir 'h%h !== 'h0", ir); end	// Vector No: 1124
assert (op === 'h00) else begin fail = 1; $display("Error 4497: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4498: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4499: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f04000:0:1:0:04:1:04000:
//------------------------

#2;
word <= 'h0000000003f04000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1126
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4500: ir 'h%h !== 'h0", ir); end	// Vector No: 1125
assert (op === 'h04) else begin fail = 1; $display("Error 4501: op 'h%h !== 'h04", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4502: extop 'h%h !== 1", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 4503: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000000003f04000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f04000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1127
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4504: ir 'h%h !== 'h0", ir); end	// Vector No: 1126
assert (op === 'h00) else begin fail = 1; $display("Error 4505: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4506: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4507: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f04000:1:1:0:03:0:00f04:
//------------------------

#2;
word <= 'h0000000003f04000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1128
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4508: ir 'h%h !== 'h0", ir); end	// Vector No: 1127
assert (op === 'h03) else begin fail = 1; $display("Error 4509: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4510: extop 'h%h !== 0", extop); end
assert (addr === 'h00f04) else begin fail = 1; $display("Error 4511: addr 'h%h !== 'h00f04", addr); end
#2;
clk <= 0;

// 03f0000000004000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000004000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1129
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4512: ir 'h%h !== 'h0", ir); end	// Vector No: 1128
assert (op === 'h00) else begin fail = 1; $display("Error 4513: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4514: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4515: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000004000:0:1:0:00:0:04000:
//------------------------

#2;
word <= 'h03f0000000004000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1130
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4516: ir 'h%h !== 'h0", ir); end	// Vector No: 1129
assert (op === 'h00) else begin fail = 1; $display("Error 4517: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4518: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 4519: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 03f0000000004000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000004000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1131
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4520: ir 'h%h !== 'h3", ir); end	// Vector No: 1130
assert (op === 'hf0) else begin fail = 1; $display("Error 4521: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4522: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4523: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000004000:1:1:0:00:0:00004:
//------------------------

#2;
word <= 'h03f0000000004000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1132
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4524: ir 'h%h !== 'h0", ir); end	// Vector No: 1131
assert (op === 'h00) else begin fail = 1; $display("Error 4525: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4526: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 4527: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000003f08000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f08000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1133
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4528: ir 'h%h !== 'h0", ir); end	// Vector No: 1132
assert (op === 'h00) else begin fail = 1; $display("Error 4529: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4530: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4531: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f08000:0:1:0:08:1:08000:
//------------------------

#2;
word <= 'h0000000003f08000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1134
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4532: ir 'h%h !== 'h0", ir); end	// Vector No: 1133
assert (op === 'h08) else begin fail = 1; $display("Error 4533: op 'h%h !== 'h08", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4534: extop 'h%h !== 1", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 4535: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000000003f08000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f08000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1135
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4536: ir 'h%h !== 'h0", ir); end	// Vector No: 1134
assert (op === 'h00) else begin fail = 1; $display("Error 4537: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4538: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4539: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f08000:1:1:0:03:0:00f08:
//------------------------

#2;
word <= 'h0000000003f08000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1136
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4540: ir 'h%h !== 'h0", ir); end	// Vector No: 1135
assert (op === 'h03) else begin fail = 1; $display("Error 4541: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4542: extop 'h%h !== 0", extop); end
assert (addr === 'h00f08) else begin fail = 1; $display("Error 4543: addr 'h%h !== 'h00f08", addr); end
#2;
clk <= 0;

// 03f0000000008000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000008000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1137
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4544: ir 'h%h !== 'h0", ir); end	// Vector No: 1136
assert (op === 'h00) else begin fail = 1; $display("Error 4545: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4546: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4547: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000008000:0:1:0:00:0:08000:
//------------------------

#2;
word <= 'h03f0000000008000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1138
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4548: ir 'h%h !== 'h0", ir); end	// Vector No: 1137
assert (op === 'h00) else begin fail = 1; $display("Error 4549: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4550: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 4551: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 03f0000000008000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000008000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1139
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4552: ir 'h%h !== 'h3", ir); end	// Vector No: 1138
assert (op === 'hf0) else begin fail = 1; $display("Error 4553: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4554: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4555: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000008000:1:1:0:00:0:00008:
//------------------------

#2;
word <= 'h03f0000000008000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1140
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4556: ir 'h%h !== 'h0", ir); end	// Vector No: 1139
assert (op === 'h00) else begin fail = 1; $display("Error 4557: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4558: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 4559: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000003f10000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f10000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1141
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4560: ir 'h%h !== 'h0", ir); end	// Vector No: 1140
assert (op === 'h00) else begin fail = 1; $display("Error 4561: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4562: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4563: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f10000:0:1:0:10:1:10000:
//------------------------

#2;
word <= 'h0000000003f10000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1142
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4564: ir 'h%h !== 'h0", ir); end	// Vector No: 1141
assert (op === 'h10) else begin fail = 1; $display("Error 4565: op 'h%h !== 'h10", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4566: extop 'h%h !== 1", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 4567: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0000000003f10000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f10000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1143
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4568: ir 'h%h !== 'h0", ir); end	// Vector No: 1142
assert (op === 'h00) else begin fail = 1; $display("Error 4569: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4570: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4571: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f10000:1:1:0:03:0:00f10:
//------------------------

#2;
word <= 'h0000000003f10000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1144
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4572: ir 'h%h !== 'h0", ir); end	// Vector No: 1143
assert (op === 'h03) else begin fail = 1; $display("Error 4573: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4574: extop 'h%h !== 0", extop); end
assert (addr === 'h00f10) else begin fail = 1; $display("Error 4575: addr 'h%h !== 'h00f10", addr); end
#2;
clk <= 0;

// 03f0000000010000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1145
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4576: ir 'h%h !== 'h0", ir); end	// Vector No: 1144
assert (op === 'h00) else begin fail = 1; $display("Error 4577: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4578: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4579: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000010000:0:1:0:00:0:10000:
//------------------------

#2;
word <= 'h03f0000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1146
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4580: ir 'h%h !== 'h0", ir); end	// Vector No: 1145
assert (op === 'h00) else begin fail = 1; $display("Error 4581: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4582: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 4583: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 03f0000000010000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1147
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4584: ir 'h%h !== 'h3", ir); end	// Vector No: 1146
assert (op === 'hf0) else begin fail = 1; $display("Error 4585: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4586: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4587: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000010000:1:1:0:00:0:00010:
//------------------------

#2;
word <= 'h03f0000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1148
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4588: ir 'h%h !== 'h0", ir); end	// Vector No: 1147
assert (op === 'h00) else begin fail = 1; $display("Error 4589: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4590: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 4591: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000000003f20000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f20000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1149
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4592: ir 'h%h !== 'h0", ir); end	// Vector No: 1148
assert (op === 'h00) else begin fail = 1; $display("Error 4593: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4594: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4595: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f20000:0:1:0:20:1:20000:
//------------------------

#2;
word <= 'h0000000003f20000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1150
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4596: ir 'h%h !== 'h0", ir); end	// Vector No: 1149
assert (op === 'h20) else begin fail = 1; $display("Error 4597: op 'h%h !== 'h20", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4598: extop 'h%h !== 1", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 4599: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0000000003f20000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f20000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1151
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4600: ir 'h%h !== 'h0", ir); end	// Vector No: 1150
assert (op === 'h00) else begin fail = 1; $display("Error 4601: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4602: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4603: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f20000:1:1:0:03:0:00f20:
//------------------------

#2;
word <= 'h0000000003f20000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1152
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4604: ir 'h%h !== 'h0", ir); end	// Vector No: 1151
assert (op === 'h03) else begin fail = 1; $display("Error 4605: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4606: extop 'h%h !== 0", extop); end
assert (addr === 'h00f20) else begin fail = 1; $display("Error 4607: addr 'h%h !== 'h00f20", addr); end
#2;
clk <= 0;

// 03f0000000020000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000020000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1153
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4608: ir 'h%h !== 'h0", ir); end	// Vector No: 1152
assert (op === 'h00) else begin fail = 1; $display("Error 4609: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4610: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4611: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000020000:0:1:0:00:0:20000:
//------------------------

#2;
word <= 'h03f0000000020000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1154
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4612: ir 'h%h !== 'h0", ir); end	// Vector No: 1153
assert (op === 'h00) else begin fail = 1; $display("Error 4613: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4614: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 4615: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 03f0000000020000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000020000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1155
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4616: ir 'h%h !== 'h3", ir); end	// Vector No: 1154
assert (op === 'hf0) else begin fail = 1; $display("Error 4617: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4618: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4619: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000020000:1:1:0:00:0:00020:
//------------------------

#2;
word <= 'h03f0000000020000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1156
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4620: ir 'h%h !== 'h0", ir); end	// Vector No: 1155
assert (op === 'h00) else begin fail = 1; $display("Error 4621: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4622: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 4623: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000000003f40000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f40000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1157
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4624: ir 'h%h !== 'h0", ir); end	// Vector No: 1156
assert (op === 'h00) else begin fail = 1; $display("Error 4625: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4626: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4627: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f40000:0:1:0:40:1:40000:
//------------------------

#2;
word <= 'h0000000003f40000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1158
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4628: ir 'h%h !== 'h0", ir); end	// Vector No: 1157
assert (op === 'h40) else begin fail = 1; $display("Error 4629: op 'h%h !== 'h40", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4630: extop 'h%h !== 1", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 4631: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0000000003f40000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f40000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1159
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4632: ir 'h%h !== 'h0", ir); end	// Vector No: 1158
assert (op === 'h00) else begin fail = 1; $display("Error 4633: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4634: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4635: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f40000:1:1:0:03:0:00f40:
//------------------------

#2;
word <= 'h0000000003f40000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1160
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4636: ir 'h%h !== 'h0", ir); end	// Vector No: 1159
assert (op === 'h03) else begin fail = 1; $display("Error 4637: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4638: extop 'h%h !== 0", extop); end
assert (addr === 'h00f40) else begin fail = 1; $display("Error 4639: addr 'h%h !== 'h00f40", addr); end
#2;
clk <= 0;

// 03f0000000040000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000040000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1161
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4640: ir 'h%h !== 'h0", ir); end	// Vector No: 1160
assert (op === 'h00) else begin fail = 1; $display("Error 4641: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4642: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4643: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000040000:0:1:0:00:0:40000:
//------------------------

#2;
word <= 'h03f0000000040000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1162
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4644: ir 'h%h !== 'h0", ir); end	// Vector No: 1161
assert (op === 'h00) else begin fail = 1; $display("Error 4645: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4646: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 4647: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 03f0000000040000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000040000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1163
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4648: ir 'h%h !== 'h3", ir); end	// Vector No: 1162
assert (op === 'hf0) else begin fail = 1; $display("Error 4649: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4650: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4651: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000040000:1:1:0:00:0:00040:
//------------------------

#2;
word <= 'h03f0000000040000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1164
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4652: ir 'h%h !== 'h0", ir); end	// Vector No: 1163
assert (op === 'h00) else begin fail = 1; $display("Error 4653: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4654: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 4655: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000000003f80000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f80000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1165
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4656: ir 'h%h !== 'h0", ir); end	// Vector No: 1164
assert (op === 'h00) else begin fail = 1; $display("Error 4657: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4658: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4659: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f80000:0:1:0:80:1:80000:
//------------------------

#2;
word <= 'h0000000003f80000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1166
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4660: ir 'h%h !== 'h0", ir); end	// Vector No: 1165
assert (op === 'h80) else begin fail = 1; $display("Error 4661: op 'h%h !== 'h80", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4662: extop 'h%h !== 1", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 4663: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0000000003f80000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f80000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1167
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4664: ir 'h%h !== 'h0", ir); end	// Vector No: 1166
assert (op === 'h00) else begin fail = 1; $display("Error 4665: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4666: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4667: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f80000:1:1:0:03:0:00f80:
//------------------------

#2;
word <= 'h0000000003f80000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1168
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4668: ir 'h%h !== 'h0", ir); end	// Vector No: 1167
assert (op === 'h03) else begin fail = 1; $display("Error 4669: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4670: extop 'h%h !== 0", extop); end
assert (addr === 'h00f80) else begin fail = 1; $display("Error 4671: addr 'h%h !== 'h00f80", addr); end
#2;
clk <= 0;

// 03f0000000080000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000080000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1169
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4672: ir 'h%h !== 'h0", ir); end	// Vector No: 1168
assert (op === 'h00) else begin fail = 1; $display("Error 4673: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4674: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4675: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000080000:0:1:0:00:0:80000:
//------------------------

#2;
word <= 'h03f0000000080000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1170
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4676: ir 'h%h !== 'h0", ir); end	// Vector No: 1169
assert (op === 'h00) else begin fail = 1; $display("Error 4677: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4678: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 4679: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 03f0000000080000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000080000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1171
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4680: ir 'h%h !== 'h3", ir); end	// Vector No: 1170
assert (op === 'hf0) else begin fail = 1; $display("Error 4681: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4682: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4683: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000080000:1:1:0:00:0:00080:
//------------------------

#2;
word <= 'h03f0000000080000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1172
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4684: ir 'h%h !== 'h0", ir); end	// Vector No: 1171
assert (op === 'h00) else begin fail = 1; $display("Error 4685: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4686: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 4687: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000000003f00000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1173
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4688: ir 'h%h !== 'h0", ir); end	// Vector No: 1172
assert (op === 'h00) else begin fail = 1; $display("Error 4689: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4690: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4691: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1174
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4692: ir 'h%h !== 'h0", ir); end	// Vector No: 1173
assert (op === 'h00) else begin fail = 1; $display("Error 4693: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4694: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4695: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1175
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4696: ir 'h%h !== 'h0", ir); end	// Vector No: 1174
assert (op === 'h00) else begin fail = 1; $display("Error 4697: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4698: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4699: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1176
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4700: ir 'h%h !== 'h0", ir); end	// Vector No: 1175
assert (op === 'h03) else begin fail = 1; $display("Error 4701: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4702: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4703: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000100000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1177
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4704: ir 'h%h !== 'h0", ir); end	// Vector No: 1176
assert (op === 'h00) else begin fail = 1; $display("Error 4705: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4706: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4707: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000100000:0:1:0:01:0:00000:
//------------------------

#2;
word <= 'h03f0000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1178
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4708: ir 'h%h !== 'h0", ir); end	// Vector No: 1177
assert (op === 'h01) else begin fail = 1; $display("Error 4709: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4710: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4711: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000100000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1179
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4712: ir 'h%h !== 'h3", ir); end	// Vector No: 1178
assert (op === 'hf0) else begin fail = 1; $display("Error 4713: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4714: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4715: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000100000:1:1:0:00:0:00100:
//------------------------

#2;
word <= 'h03f0000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1180
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4716: ir 'h%h !== 'h0", ir); end	// Vector No: 1179
assert (op === 'h00) else begin fail = 1; $display("Error 4717: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4718: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 4719: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 03f0000000200000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000200000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1181
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4720: ir 'h%h !== 'h0", ir); end	// Vector No: 1180
assert (op === 'h00) else begin fail = 1; $display("Error 4721: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4722: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4723: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000200000:0:1:0:02:0:00000:
//------------------------

#2;
word <= 'h03f0000000200000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1182
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4724: ir 'h%h !== 'h0", ir); end	// Vector No: 1181
assert (op === 'h02) else begin fail = 1; $display("Error 4725: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4726: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4727: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000200000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000200000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1183
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4728: ir 'h%h !== 'h3", ir); end	// Vector No: 1182
assert (op === 'hf0) else begin fail = 1; $display("Error 4729: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4730: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4731: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000200000:1:1:0:00:0:00200:
//------------------------

#2;
word <= 'h03f0000000200000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1184
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4732: ir 'h%h !== 'h0", ir); end	// Vector No: 1183
assert (op === 'h00) else begin fail = 1; $display("Error 4733: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4734: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 4735: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 03f0000000400000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000400000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1185
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4736: ir 'h%h !== 'h0", ir); end	// Vector No: 1184
assert (op === 'h00) else begin fail = 1; $display("Error 4737: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4738: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4739: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000400000:0:1:0:04:0:00000:
//------------------------

#2;
word <= 'h03f0000000400000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1186
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4740: ir 'h%h !== 'h0", ir); end	// Vector No: 1185
assert (op === 'h04) else begin fail = 1; $display("Error 4741: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4742: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4743: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000400000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000400000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1187
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4744: ir 'h%h !== 'h3", ir); end	// Vector No: 1186
assert (op === 'hf0) else begin fail = 1; $display("Error 4745: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4746: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4747: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000400000:1:1:0:00:0:00400:
//------------------------

#2;
word <= 'h03f0000000400000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1188
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4748: ir 'h%h !== 'h0", ir); end	// Vector No: 1187
assert (op === 'h00) else begin fail = 1; $display("Error 4749: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4750: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 4751: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 03f0000000800000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000800000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1189
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4752: ir 'h%h !== 'h0", ir); end	// Vector No: 1188
assert (op === 'h00) else begin fail = 1; $display("Error 4753: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4754: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4755: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000800000:0:1:0:08:0:00000:
//------------------------

#2;
word <= 'h03f0000000800000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1190
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4756: ir 'h%h !== 'h0", ir); end	// Vector No: 1189
assert (op === 'h08) else begin fail = 1; $display("Error 4757: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4758: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4759: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000800000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000800000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1191
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4760: ir 'h%h !== 'h3", ir); end	// Vector No: 1190
assert (op === 'hf0) else begin fail = 1; $display("Error 4761: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4762: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4763: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000800000:1:1:0:00:0:00800:
//------------------------

#2;
word <= 'h03f0000000800000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1192
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4764: ir 'h%h !== 'h0", ir); end	// Vector No: 1191
assert (op === 'h00) else begin fail = 1; $display("Error 4765: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4766: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 4767: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 03f0000001000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1193
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4768: ir 'h%h !== 'h0", ir); end	// Vector No: 1192
assert (op === 'h00) else begin fail = 1; $display("Error 4769: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4770: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4771: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000001000000:0:1:0:10:0:00000:
//------------------------

#2;
word <= 'h03f0000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1194
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4772: ir 'h%h !== 'h0", ir); end	// Vector No: 1193
assert (op === 'h10) else begin fail = 1; $display("Error 4773: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4774: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4775: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000001000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1195
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4776: ir 'h%h !== 'h3", ir); end	// Vector No: 1194
assert (op === 'hf0) else begin fail = 1; $display("Error 4777: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4778: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4779: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000001000000:1:1:0:01:0:00000:
//------------------------

#2;
word <= 'h03f0000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1196
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4780: ir 'h%h !== 'h0", ir); end	// Vector No: 1195
assert (op === 'h01) else begin fail = 1; $display("Error 4781: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4782: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4783: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000002000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000002000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1197
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4784: ir 'h%h !== 'h0", ir); end	// Vector No: 1196
assert (op === 'h00) else begin fail = 1; $display("Error 4785: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4786: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4787: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000002000000:0:1:0:20:0:00000:
//------------------------

#2;
word <= 'h03f0000002000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1198
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4788: ir 'h%h !== 'h0", ir); end	// Vector No: 1197
assert (op === 'h20) else begin fail = 1; $display("Error 4789: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4790: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4791: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000002000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000002000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1199
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4792: ir 'h%h !== 'h3", ir); end	// Vector No: 1198
assert (op === 'hf0) else begin fail = 1; $display("Error 4793: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4794: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4795: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000002000000:1:1:0:02:0:00000:
//------------------------

#2;
word <= 'h03f0000002000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1200
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4796: ir 'h%h !== 'h0", ir); end	// Vector No: 1199
assert (op === 'h02) else begin fail = 1; $display("Error 4797: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4798: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4799: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000004000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000004000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1201
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4800: ir 'h%h !== 'h0", ir); end	// Vector No: 1200
assert (op === 'h00) else begin fail = 1; $display("Error 4801: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4802: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4803: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000004000000:0:1:0:40:0:00000:
//------------------------

#2;
word <= 'h03f0000004000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1202
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4804: ir 'h%h !== 'h0", ir); end	// Vector No: 1201
assert (op === 'h40) else begin fail = 1; $display("Error 4805: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4806: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4807: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000004000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000004000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1203
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4808: ir 'h%h !== 'h3", ir); end	// Vector No: 1202
assert (op === 'hf0) else begin fail = 1; $display("Error 4809: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4810: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4811: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000004000000:1:1:0:04:0:00000:
//------------------------

#2;
word <= 'h03f0000004000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1204
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4812: ir 'h%h !== 'h0", ir); end	// Vector No: 1203
assert (op === 'h04) else begin fail = 1; $display("Error 4813: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4814: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4815: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000008000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000008000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1205
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4816: ir 'h%h !== 'h0", ir); end	// Vector No: 1204
assert (op === 'h00) else begin fail = 1; $display("Error 4817: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4818: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4819: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000008000000:0:1:0:80:0:00000:
//------------------------

#2;
word <= 'h03f0000008000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1206
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4820: ir 'h%h !== 'h0", ir); end	// Vector No: 1205
assert (op === 'h80) else begin fail = 1; $display("Error 4821: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4822: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4823: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000008000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000008000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1207
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4824: ir 'h%h !== 'h3", ir); end	// Vector No: 1206
assert (op === 'hf0) else begin fail = 1; $display("Error 4825: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4826: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4827: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000008000000:1:1:0:08:0:00000:
//------------------------

#2;
word <= 'h03f0000008000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1208
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4828: ir 'h%h !== 'h0", ir); end	// Vector No: 1207
assert (op === 'h08) else begin fail = 1; $display("Error 4829: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4830: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4831: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000013f00000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000013f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1209
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4832: ir 'h%h !== 'h0", ir); end	// Vector No: 1208
assert (op === 'h00) else begin fail = 1; $display("Error 4833: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4834: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4835: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000013f00000:0:1:1:00:1:00000:
//------------------------

#2;
word <= 'h0000000013f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1210
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 4836: ir 'h%h !== 'h1", ir); end	// Vector No: 1209
assert (op === 'h00) else begin fail = 1; $display("Error 4837: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4838: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4839: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000013f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000013f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1211
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4840: ir 'h%h !== 'h0", ir); end	// Vector No: 1210
assert (op === 'h00) else begin fail = 1; $display("Error 4841: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4842: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4843: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000013f00000:1:1:0:13:0:00f00:
//------------------------

#2;
word <= 'h0000000013f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1212
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4844: ir 'h%h !== 'h0", ir); end	// Vector No: 1211
assert (op === 'h13) else begin fail = 1; $display("Error 4845: op 'h%h !== 'h13", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4846: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4847: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000010000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1213
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4848: ir 'h%h !== 'h0", ir); end	// Vector No: 1212
assert (op === 'h00) else begin fail = 1; $display("Error 4849: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4850: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4851: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000010000000:0:1:1:00:0:00000:
//------------------------

#2;
word <= 'h03f0000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1214
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 4852: ir 'h%h !== 'h1", ir); end	// Vector No: 1213
assert (op === 'h00) else begin fail = 1; $display("Error 4853: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4854: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4855: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000010000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1215
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4856: ir 'h%h !== 'h3", ir); end	// Vector No: 1214
assert (op === 'hf0) else begin fail = 1; $display("Error 4857: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4858: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4859: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000010000000:1:1:0:10:0:00000:
//------------------------

#2;
word <= 'h03f0000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1216
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4860: ir 'h%h !== 'h0", ir); end	// Vector No: 1215
assert (op === 'h10) else begin fail = 1; $display("Error 4861: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4862: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4863: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000023f00000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000023f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1217
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4864: ir 'h%h !== 'h0", ir); end	// Vector No: 1216
assert (op === 'h00) else begin fail = 1; $display("Error 4865: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4866: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4867: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000023f00000:0:1:2:00:1:00000:
//------------------------

#2;
word <= 'h0000000023f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1218
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 4868: ir 'h%h !== 'h2", ir); end	// Vector No: 1217
assert (op === 'h00) else begin fail = 1; $display("Error 4869: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4870: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4871: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000023f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000023f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1219
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4872: ir 'h%h !== 'h0", ir); end	// Vector No: 1218
assert (op === 'h00) else begin fail = 1; $display("Error 4873: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4874: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4875: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000023f00000:1:1:0:23:0:00f00:
//------------------------

#2;
word <= 'h0000000023f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1220
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4876: ir 'h%h !== 'h0", ir); end	// Vector No: 1219
assert (op === 'h23) else begin fail = 1; $display("Error 4877: op 'h%h !== 'h23", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4878: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4879: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000020000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000020000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1221
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4880: ir 'h%h !== 'h0", ir); end	// Vector No: 1220
assert (op === 'h00) else begin fail = 1; $display("Error 4881: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4882: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4883: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000020000000:0:1:2:00:0:00000:
//------------------------

#2;
word <= 'h03f0000020000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1222
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 4884: ir 'h%h !== 'h2", ir); end	// Vector No: 1221
assert (op === 'h00) else begin fail = 1; $display("Error 4885: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4886: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4887: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000020000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000020000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1223
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4888: ir 'h%h !== 'h3", ir); end	// Vector No: 1222
assert (op === 'hf0) else begin fail = 1; $display("Error 4889: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4890: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4891: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000020000000:1:1:0:20:0:00000:
//------------------------

#2;
word <= 'h03f0000020000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1224
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4892: ir 'h%h !== 'h0", ir); end	// Vector No: 1223
assert (op === 'h20) else begin fail = 1; $display("Error 4893: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4894: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4895: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000043f00000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000043f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1225
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4896: ir 'h%h !== 'h0", ir); end	// Vector No: 1224
assert (op === 'h00) else begin fail = 1; $display("Error 4897: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4898: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4899: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000043f00000:0:1:4:00:1:00000:
//------------------------

#2;
word <= 'h0000000043f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1226
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 4900: ir 'h%h !== 'h4", ir); end	// Vector No: 1225
assert (op === 'h00) else begin fail = 1; $display("Error 4901: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4902: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4903: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000043f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000043f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1227
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4904: ir 'h%h !== 'h0", ir); end	// Vector No: 1226
assert (op === 'h00) else begin fail = 1; $display("Error 4905: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4906: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4907: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000043f00000:1:1:0:43:0:07f00:
//------------------------

#2;
word <= 'h0000000043f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1228
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4908: ir 'h%h !== 'h0", ir); end	// Vector No: 1227
assert (op === 'h43) else begin fail = 1; $display("Error 4909: op 'h%h !== 'h43", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4910: extop 'h%h !== 0", extop); end
assert (addr === 'h07f00) else begin fail = 1; $display("Error 4911: addr 'h%h !== 'h07f00", addr); end
#2;
clk <= 0;

// 03f0000040000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000040000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1229
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4912: ir 'h%h !== 'h0", ir); end	// Vector No: 1228
assert (op === 'h00) else begin fail = 1; $display("Error 4913: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4914: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4915: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000040000000:0:1:4:00:0:00000:
//------------------------

#2;
word <= 'h03f0000040000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1230
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 4916: ir 'h%h !== 'h4", ir); end	// Vector No: 1229
assert (op === 'h00) else begin fail = 1; $display("Error 4917: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4918: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4919: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000040000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000040000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1231
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4920: ir 'h%h !== 'h3", ir); end	// Vector No: 1230
assert (op === 'hf0) else begin fail = 1; $display("Error 4921: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4922: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4923: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000040000000:1:1:0:40:0:07000:
//------------------------

#2;
word <= 'h03f0000040000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1232
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4924: ir 'h%h !== 'h0", ir); end	// Vector No: 1231
assert (op === 'h40) else begin fail = 1; $display("Error 4925: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4926: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 4927: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0000000083f00000:0:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000083f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1233
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4928: ir 'h%h !== 'h0", ir); end	// Vector No: 1232
assert (op === 'h00) else begin fail = 1; $display("Error 4929: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4930: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4931: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000083f00000:0:1:8:00:1:00000:
//------------------------

#2;
word <= 'h0000000083f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1234
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 4932: ir 'h%h !== 'h8", ir); end	// Vector No: 1233
assert (op === 'h00) else begin fail = 1; $display("Error 4933: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4934: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4935: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000083f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000083f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1235
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4936: ir 'h%h !== 'h0", ir); end	// Vector No: 1234
assert (op === 'h00) else begin fail = 1; $display("Error 4937: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4938: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4939: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000083f00000:1:1:0:80:0:03f00:
//------------------------

#2;
word <= 'h0000000083f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1236
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4940: ir 'h%h !== 'h0", ir); end	// Vector No: 1235
assert (op === 'h80) else begin fail = 1; $display("Error 4941: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4942: extop 'h%h !== 0", extop); end
assert (addr === 'h03f00) else begin fail = 1; $display("Error 4943: addr 'h%h !== 'h03f00", addr); end
#2;
clk <= 0;

// 03f0000080000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000080000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1237
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4944: ir 'h%h !== 'h0", ir); end	// Vector No: 1236
assert (op === 'h00) else begin fail = 1; $display("Error 4945: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4946: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4947: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000080000000:0:1:8:00:0:00000:
//------------------------

#2;
word <= 'h03f0000080000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1238
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 4948: ir 'h%h !== 'h8", ir); end	// Vector No: 1237
assert (op === 'h00) else begin fail = 1; $display("Error 4949: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4950: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4951: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000080000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000080000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1239
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4952: ir 'h%h !== 'h3", ir); end	// Vector No: 1238
assert (op === 'hf0) else begin fail = 1; $display("Error 4953: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4954: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4955: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000080000000:1:1:0:80:0:00000:
//------------------------

#2;
word <= 'h03f0000080000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1240
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4956: ir 'h%h !== 'h0", ir); end	// Vector No: 1239
assert (op === 'h80) else begin fail = 1; $display("Error 4957: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4958: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4959: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000103f00000:0:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000000103f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1241
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4960: ir 'h%h !== 'h0", ir); end	// Vector No: 1240
assert (op === 'h00) else begin fail = 1; $display("Error 4961: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4962: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 4963: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000000103f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000000103f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1242
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4964: ir 'h%h !== 'h0", ir); end	// Vector No: 1241
assert (op === 'h00) else begin fail = 1; $display("Error 4965: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4966: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4967: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000103f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000103f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1243
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4968: ir 'h%h !== 'h0", ir); end	// Vector No: 1242
assert (op === 'h00) else begin fail = 1; $display("Error 4969: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4970: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4971: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000103f00000:1:1:1:03:0:00f00:
//------------------------

#2;
word <= 'h0000000103f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1244
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 4972: ir 'h%h !== 'h1", ir); end	// Vector No: 1243
assert (op === 'h03) else begin fail = 1; $display("Error 4973: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4974: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 4975: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000100000000:0:0:0:00:1:00001:
//------------------------

#2;
word <= 'h03f0000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1245
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4976: ir 'h%h !== 'h0", ir); end	// Vector No: 1244
assert (op === 'h00) else begin fail = 1; $display("Error 4977: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4978: extop 'h%h !== 1", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 4979: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 03f0000100000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1246
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4980: ir 'h%h !== 'h0", ir); end	// Vector No: 1245
assert (op === 'h00) else begin fail = 1; $display("Error 4981: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4982: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4983: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000100000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1247
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 4984: ir 'h%h !== 'h3", ir); end	// Vector No: 1246
assert (op === 'hf0) else begin fail = 1; $display("Error 4985: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4986: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4987: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000100000000:1:1:1:00:0:00000:
//------------------------

#2;
word <= 'h03f0000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1248
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 4988: ir 'h%h !== 'h1", ir); end	// Vector No: 1247
assert (op === 'h00) else begin fail = 1; $display("Error 4989: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4990: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4991: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000203f00000:0:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000000203f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1249
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4992: ir 'h%h !== 'h0", ir); end	// Vector No: 1248
assert (op === 'h00) else begin fail = 1; $display("Error 4993: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 4994: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 4995: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000000203f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000000203f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1250
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 4996: ir 'h%h !== 'h0", ir); end	// Vector No: 1249
assert (op === 'h00) else begin fail = 1; $display("Error 4997: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 4998: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 4999: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000203f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000203f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1251
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5000: ir 'h%h !== 'h0", ir); end	// Vector No: 1250
assert (op === 'h00) else begin fail = 1; $display("Error 5001: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5002: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5003: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000203f00000:1:1:2:03:0:00f00:
//------------------------

#2;
word <= 'h0000000203f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1252
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 5004: ir 'h%h !== 'h2", ir); end	// Vector No: 1251
assert (op === 'h03) else begin fail = 1; $display("Error 5005: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5006: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5007: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000200000000:0:0:0:00:1:00002:
//------------------------

#2;
word <= 'h03f0000200000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1253
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5008: ir 'h%h !== 'h0", ir); end	// Vector No: 1252
assert (op === 'h00) else begin fail = 1; $display("Error 5009: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5010: extop 'h%h !== 1", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 5011: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 03f0000200000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000200000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1254
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5012: ir 'h%h !== 'h0", ir); end	// Vector No: 1253
assert (op === 'h00) else begin fail = 1; $display("Error 5013: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5014: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5015: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000200000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000200000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1255
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5016: ir 'h%h !== 'h3", ir); end	// Vector No: 1254
assert (op === 'hf0) else begin fail = 1; $display("Error 5017: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5018: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5019: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000200000000:1:1:2:00:0:00000:
//------------------------

#2;
word <= 'h03f0000200000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1256
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 5020: ir 'h%h !== 'h2", ir); end	// Vector No: 1255
assert (op === 'h00) else begin fail = 1; $display("Error 5021: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5022: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5023: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000403f00000:0:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000000403f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1257
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5024: ir 'h%h !== 'h0", ir); end	// Vector No: 1256
assert (op === 'h00) else begin fail = 1; $display("Error 5025: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5026: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 5027: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000000403f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000000403f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1258
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5028: ir 'h%h !== 'h0", ir); end	// Vector No: 1257
assert (op === 'h00) else begin fail = 1; $display("Error 5029: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5030: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5031: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000403f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000403f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1259
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5032: ir 'h%h !== 'h0", ir); end	// Vector No: 1258
assert (op === 'h00) else begin fail = 1; $display("Error 5033: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5034: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5035: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000403f00000:1:1:4:03:0:00f00:
//------------------------

#2;
word <= 'h0000000403f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1260
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 5036: ir 'h%h !== 'h4", ir); end	// Vector No: 1259
assert (op === 'h03) else begin fail = 1; $display("Error 5037: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5038: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5039: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000400000000:0:0:0:00:1:00004:
//------------------------

#2;
word <= 'h03f0000400000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1261
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5040: ir 'h%h !== 'h0", ir); end	// Vector No: 1260
assert (op === 'h00) else begin fail = 1; $display("Error 5041: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5042: extop 'h%h !== 1", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 5043: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 03f0000400000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000400000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1262
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5044: ir 'h%h !== 'h0", ir); end	// Vector No: 1261
assert (op === 'h00) else begin fail = 1; $display("Error 5045: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5046: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5047: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000400000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000400000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1263
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5048: ir 'h%h !== 'h3", ir); end	// Vector No: 1262
assert (op === 'hf0) else begin fail = 1; $display("Error 5049: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5050: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5051: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000400000000:1:1:4:00:0:00000:
//------------------------

#2;
word <= 'h03f0000400000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1264
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 5052: ir 'h%h !== 'h4", ir); end	// Vector No: 1263
assert (op === 'h00) else begin fail = 1; $display("Error 5053: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5054: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5055: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000803f00000:0:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000000803f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1265
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5056: ir 'h%h !== 'h0", ir); end	// Vector No: 1264
assert (op === 'h00) else begin fail = 1; $display("Error 5057: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5058: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 5059: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000000803f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000000803f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1266
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5060: ir 'h%h !== 'h0", ir); end	// Vector No: 1265
assert (op === 'h00) else begin fail = 1; $display("Error 5061: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5062: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5063: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000803f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0000000803f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1267
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5064: ir 'h%h !== 'h0", ir); end	// Vector No: 1266
assert (op === 'h00) else begin fail = 1; $display("Error 5065: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5066: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5067: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000000803f00000:1:1:8:03:0:00f00:
//------------------------

#2;
word <= 'h0000000803f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1268
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 5068: ir 'h%h !== 'h8", ir); end	// Vector No: 1267
assert (op === 'h03) else begin fail = 1; $display("Error 5069: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5070: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5071: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000800000000:0:0:0:00:1:00008:
//------------------------

#2;
word <= 'h03f0000800000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1269
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5072: ir 'h%h !== 'h0", ir); end	// Vector No: 1268
assert (op === 'h00) else begin fail = 1; $display("Error 5073: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5074: extop 'h%h !== 1", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 5075: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 03f0000800000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000800000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1270
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5076: ir 'h%h !== 'h0", ir); end	// Vector No: 1269
assert (op === 'h00) else begin fail = 1; $display("Error 5077: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5078: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5079: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000800000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000800000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1271
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5080: ir 'h%h !== 'h3", ir); end	// Vector No: 1270
assert (op === 'hf0) else begin fail = 1; $display("Error 5081: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5082: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5083: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000800000000:1:1:8:00:0:00000:
//------------------------

#2;
word <= 'h03f0000800000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1272
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 5084: ir 'h%h !== 'h8", ir); end	// Vector No: 1271
assert (op === 'h00) else begin fail = 1; $display("Error 5085: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5086: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5087: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001003f00000:0:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000001003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1273
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5088: ir 'h%h !== 'h0", ir); end	// Vector No: 1272
assert (op === 'h00) else begin fail = 1; $display("Error 5089: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5090: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 5091: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000001003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000001003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1274
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5092: ir 'h%h !== 'h0", ir); end	// Vector No: 1273
assert (op === 'h00) else begin fail = 1; $display("Error 5093: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5094: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5095: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000001003f00000:1:0:0:00:0:00001:
//------------------------

#2;
word <= 'h0000001003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1275
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5096: ir 'h%h !== 'h0", ir); end	// Vector No: 1274
assert (op === 'h00) else begin fail = 1; $display("Error 5097: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5098: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 5099: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 0000001003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000001003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1276
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5100: ir 'h%h !== 'h0", ir); end	// Vector No: 1275
assert (op === 'h03) else begin fail = 1; $display("Error 5101: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5102: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5103: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0001000000000:0:0:0:00:1:00010:
//------------------------

#2;
word <= 'h03f0001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1277
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5104: ir 'h%h !== 'h0", ir); end	// Vector No: 1276
assert (op === 'h00) else begin fail = 1; $display("Error 5105: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5106: extop 'h%h !== 1", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 5107: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 03f0001000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1278
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5108: ir 'h%h !== 'h0", ir); end	// Vector No: 1277
assert (op === 'h00) else begin fail = 1; $display("Error 5109: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5110: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5111: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0001000000000:1:0:3:f0:0:00001:
//------------------------

#2;
word <= 'h03f0001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1279
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5112: ir 'h%h !== 'h3", ir); end	// Vector No: 1278
assert (op === 'hf0) else begin fail = 1; $display("Error 5113: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5114: extop 'h%h !== 0", extop); end
assert (addr === 'h00001) else begin fail = 1; $display("Error 5115: addr 'h%h !== 'h00001", addr); end
#2;
clk <= 0;

// 03f0001000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1280
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5116: ir 'h%h !== 'h0", ir); end	// Vector No: 1279
assert (op === 'h00) else begin fail = 1; $display("Error 5117: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5118: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5119: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002003f00000:0:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000002003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1281
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5120: ir 'h%h !== 'h0", ir); end	// Vector No: 1280
assert (op === 'h00) else begin fail = 1; $display("Error 5121: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5122: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 5123: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000002003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000002003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1282
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5124: ir 'h%h !== 'h0", ir); end	// Vector No: 1281
assert (op === 'h00) else begin fail = 1; $display("Error 5125: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5126: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5127: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000002003f00000:1:0:0:00:0:00002:
//------------------------

#2;
word <= 'h0000002003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1283
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5128: ir 'h%h !== 'h0", ir); end	// Vector No: 1282
assert (op === 'h00) else begin fail = 1; $display("Error 5129: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5130: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 5131: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 0000002003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000002003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1284
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5132: ir 'h%h !== 'h0", ir); end	// Vector No: 1283
assert (op === 'h03) else begin fail = 1; $display("Error 5133: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5134: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5135: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0002000000000:0:0:0:00:1:00020:
//------------------------

#2;
word <= 'h03f0002000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1285
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5136: ir 'h%h !== 'h0", ir); end	// Vector No: 1284
assert (op === 'h00) else begin fail = 1; $display("Error 5137: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5138: extop 'h%h !== 1", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 5139: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 03f0002000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0002000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1286
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5140: ir 'h%h !== 'h0", ir); end	// Vector No: 1285
assert (op === 'h00) else begin fail = 1; $display("Error 5141: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5142: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5143: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0002000000000:1:0:3:f0:0:00002:
//------------------------

#2;
word <= 'h03f0002000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1287
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5144: ir 'h%h !== 'h3", ir); end	// Vector No: 1286
assert (op === 'hf0) else begin fail = 1; $display("Error 5145: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5146: extop 'h%h !== 0", extop); end
assert (addr === 'h00002) else begin fail = 1; $display("Error 5147: addr 'h%h !== 'h00002", addr); end
#2;
clk <= 0;

// 03f0002000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0002000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1288
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5148: ir 'h%h !== 'h0", ir); end	// Vector No: 1287
assert (op === 'h00) else begin fail = 1; $display("Error 5149: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5150: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5151: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004003f00000:0:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000004003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1289
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5152: ir 'h%h !== 'h0", ir); end	// Vector No: 1288
assert (op === 'h00) else begin fail = 1; $display("Error 5153: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5154: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 5155: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000004003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000004003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1290
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5156: ir 'h%h !== 'h0", ir); end	// Vector No: 1289
assert (op === 'h00) else begin fail = 1; $display("Error 5157: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5158: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5159: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000004003f00000:1:0:0:00:0:00004:
//------------------------

#2;
word <= 'h0000004003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1291
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5160: ir 'h%h !== 'h0", ir); end	// Vector No: 1290
assert (op === 'h00) else begin fail = 1; $display("Error 5161: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5162: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 5163: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 0000004003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000004003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1292
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5164: ir 'h%h !== 'h0", ir); end	// Vector No: 1291
assert (op === 'h03) else begin fail = 1; $display("Error 5165: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5166: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5167: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0004000000000:0:0:0:00:1:00040:
//------------------------

#2;
word <= 'h03f0004000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1293
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5168: ir 'h%h !== 'h0", ir); end	// Vector No: 1292
assert (op === 'h00) else begin fail = 1; $display("Error 5169: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5170: extop 'h%h !== 1", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 5171: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 03f0004000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0004000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1294
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5172: ir 'h%h !== 'h0", ir); end	// Vector No: 1293
assert (op === 'h00) else begin fail = 1; $display("Error 5173: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5174: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5175: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0004000000000:1:0:3:f0:0:00004:
//------------------------

#2;
word <= 'h03f0004000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1295
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5176: ir 'h%h !== 'h3", ir); end	// Vector No: 1294
assert (op === 'hf0) else begin fail = 1; $display("Error 5177: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5178: extop 'h%h !== 0", extop); end
assert (addr === 'h00004) else begin fail = 1; $display("Error 5179: addr 'h%h !== 'h00004", addr); end
#2;
clk <= 0;

// 03f0004000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0004000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1296
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5180: ir 'h%h !== 'h0", ir); end	// Vector No: 1295
assert (op === 'h00) else begin fail = 1; $display("Error 5181: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5182: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5183: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008003f00000:0:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000008003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1297
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5184: ir 'h%h !== 'h0", ir); end	// Vector No: 1296
assert (op === 'h00) else begin fail = 1; $display("Error 5185: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5186: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 5187: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000008003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000008003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1298
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5188: ir 'h%h !== 'h0", ir); end	// Vector No: 1297
assert (op === 'h00) else begin fail = 1; $display("Error 5189: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5190: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5191: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000008003f00000:1:0:0:00:0:00008:
//------------------------

#2;
word <= 'h0000008003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1299
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5192: ir 'h%h !== 'h0", ir); end	// Vector No: 1298
assert (op === 'h00) else begin fail = 1; $display("Error 5193: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5194: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 5195: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 0000008003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000008003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1300
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5196: ir 'h%h !== 'h0", ir); end	// Vector No: 1299
assert (op === 'h03) else begin fail = 1; $display("Error 5197: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5198: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5199: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0008000000000:0:0:0:00:1:00080:
//------------------------

#2;
word <= 'h03f0008000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1301
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5200: ir 'h%h !== 'h0", ir); end	// Vector No: 1300
assert (op === 'h00) else begin fail = 1; $display("Error 5201: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5202: extop 'h%h !== 1", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 5203: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 03f0008000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0008000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1302
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5204: ir 'h%h !== 'h0", ir); end	// Vector No: 1301
assert (op === 'h00) else begin fail = 1; $display("Error 5205: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5206: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5207: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0008000000000:1:0:3:f0:0:00008:
//------------------------

#2;
word <= 'h03f0008000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1303
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5208: ir 'h%h !== 'h3", ir); end	// Vector No: 1302
assert (op === 'hf0) else begin fail = 1; $display("Error 5209: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5210: extop 'h%h !== 0", extop); end
assert (addr === 'h00008) else begin fail = 1; $display("Error 5211: addr 'h%h !== 'h00008", addr); end
#2;
clk <= 0;

// 03f0008000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0008000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1304
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5212: ir 'h%h !== 'h0", ir); end	// Vector No: 1303
assert (op === 'h00) else begin fail = 1; $display("Error 5213: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5214: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5215: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010003f00000:0:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000010003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1305
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5216: ir 'h%h !== 'h0", ir); end	// Vector No: 1304
assert (op === 'h00) else begin fail = 1; $display("Error 5217: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5218: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 5219: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000010003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000010003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1306
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5220: ir 'h%h !== 'h0", ir); end	// Vector No: 1305
assert (op === 'h00) else begin fail = 1; $display("Error 5221: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5222: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5223: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000010003f00000:1:0:0:00:0:00010:
//------------------------

#2;
word <= 'h0000010003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1307
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5224: ir 'h%h !== 'h0", ir); end	// Vector No: 1306
assert (op === 'h00) else begin fail = 1; $display("Error 5225: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5226: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 5227: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 0000010003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000010003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1308
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5228: ir 'h%h !== 'h0", ir); end	// Vector No: 1307
assert (op === 'h03) else begin fail = 1; $display("Error 5229: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5230: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5231: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0010000000000:0:0:0:00:1:00100:
//------------------------

#2;
word <= 'h03f0010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1309
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5232: ir 'h%h !== 'h0", ir); end	// Vector No: 1308
assert (op === 'h00) else begin fail = 1; $display("Error 5233: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5234: extop 'h%h !== 1", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 5235: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 03f0010000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1310
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5236: ir 'h%h !== 'h0", ir); end	// Vector No: 1309
assert (op === 'h00) else begin fail = 1; $display("Error 5237: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5238: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5239: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0010000000000:1:0:3:f0:0:00010:
//------------------------

#2;
word <= 'h03f0010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1311
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5240: ir 'h%h !== 'h3", ir); end	// Vector No: 1310
assert (op === 'hf0) else begin fail = 1; $display("Error 5241: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5242: extop 'h%h !== 0", extop); end
assert (addr === 'h00010) else begin fail = 1; $display("Error 5243: addr 'h%h !== 'h00010", addr); end
#2;
clk <= 0;

// 03f0010000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1312
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5244: ir 'h%h !== 'h0", ir); end	// Vector No: 1311
assert (op === 'h00) else begin fail = 1; $display("Error 5245: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5246: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5247: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020003f00000:0:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000020003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1313
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5248: ir 'h%h !== 'h0", ir); end	// Vector No: 1312
assert (op === 'h00) else begin fail = 1; $display("Error 5249: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5250: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 5251: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000020003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000020003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1314
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5252: ir 'h%h !== 'h0", ir); end	// Vector No: 1313
assert (op === 'h00) else begin fail = 1; $display("Error 5253: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5254: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5255: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000020003f00000:1:0:0:00:0:00020:
//------------------------

#2;
word <= 'h0000020003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1315
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5256: ir 'h%h !== 'h0", ir); end	// Vector No: 1314
assert (op === 'h00) else begin fail = 1; $display("Error 5257: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5258: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 5259: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 0000020003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000020003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1316
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5260: ir 'h%h !== 'h0", ir); end	// Vector No: 1315
assert (op === 'h03) else begin fail = 1; $display("Error 5261: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5262: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5263: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0020000000000:0:0:0:00:1:00200:
//------------------------

#2;
word <= 'h03f0020000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1317
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5264: ir 'h%h !== 'h0", ir); end	// Vector No: 1316
assert (op === 'h00) else begin fail = 1; $display("Error 5265: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5266: extop 'h%h !== 1", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 5267: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 03f0020000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0020000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1318
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5268: ir 'h%h !== 'h0", ir); end	// Vector No: 1317
assert (op === 'h00) else begin fail = 1; $display("Error 5269: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5270: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5271: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0020000000000:1:0:3:f0:0:00020:
//------------------------

#2;
word <= 'h03f0020000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1319
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5272: ir 'h%h !== 'h3", ir); end	// Vector No: 1318
assert (op === 'hf0) else begin fail = 1; $display("Error 5273: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5274: extop 'h%h !== 0", extop); end
assert (addr === 'h00020) else begin fail = 1; $display("Error 5275: addr 'h%h !== 'h00020", addr); end
#2;
clk <= 0;

// 03f0020000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0020000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1320
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5276: ir 'h%h !== 'h0", ir); end	// Vector No: 1319
assert (op === 'h00) else begin fail = 1; $display("Error 5277: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5278: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5279: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040003f00000:0:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000040003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1321
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5280: ir 'h%h !== 'h0", ir); end	// Vector No: 1320
assert (op === 'h00) else begin fail = 1; $display("Error 5281: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5282: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 5283: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000040003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000040003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1322
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5284: ir 'h%h !== 'h0", ir); end	// Vector No: 1321
assert (op === 'h00) else begin fail = 1; $display("Error 5285: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5286: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5287: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000040003f00000:1:0:0:00:0:00040:
//------------------------

#2;
word <= 'h0000040003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1323
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5288: ir 'h%h !== 'h0", ir); end	// Vector No: 1322
assert (op === 'h00) else begin fail = 1; $display("Error 5289: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5290: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 5291: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 0000040003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000040003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1324
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5292: ir 'h%h !== 'h0", ir); end	// Vector No: 1323
assert (op === 'h03) else begin fail = 1; $display("Error 5293: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5294: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5295: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0040000000000:0:0:0:00:1:00400:
//------------------------

#2;
word <= 'h03f0040000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1325
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5296: ir 'h%h !== 'h0", ir); end	// Vector No: 1324
assert (op === 'h00) else begin fail = 1; $display("Error 5297: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5298: extop 'h%h !== 1", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 5299: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 03f0040000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0040000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1326
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5300: ir 'h%h !== 'h0", ir); end	// Vector No: 1325
assert (op === 'h00) else begin fail = 1; $display("Error 5301: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5302: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5303: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0040000000000:1:0:3:f0:0:00040:
//------------------------

#2;
word <= 'h03f0040000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1327
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5304: ir 'h%h !== 'h3", ir); end	// Vector No: 1326
assert (op === 'hf0) else begin fail = 1; $display("Error 5305: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5306: extop 'h%h !== 0", extop); end
assert (addr === 'h00040) else begin fail = 1; $display("Error 5307: addr 'h%h !== 'h00040", addr); end
#2;
clk <= 0;

// 03f0040000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0040000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1328
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5308: ir 'h%h !== 'h0", ir); end	// Vector No: 1327
assert (op === 'h00) else begin fail = 1; $display("Error 5309: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5310: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5311: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080003f00000:0:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000080003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1329
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5312: ir 'h%h !== 'h0", ir); end	// Vector No: 1328
assert (op === 'h00) else begin fail = 1; $display("Error 5313: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5314: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 5315: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000080003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000080003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1330
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5316: ir 'h%h !== 'h0", ir); end	// Vector No: 1329
assert (op === 'h00) else begin fail = 1; $display("Error 5317: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5318: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5319: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000080003f00000:1:0:0:00:0:00080:
//------------------------

#2;
word <= 'h0000080003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1331
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5320: ir 'h%h !== 'h0", ir); end	// Vector No: 1330
assert (op === 'h00) else begin fail = 1; $display("Error 5321: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5322: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 5323: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 0000080003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000080003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1332
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5324: ir 'h%h !== 'h0", ir); end	// Vector No: 1331
assert (op === 'h03) else begin fail = 1; $display("Error 5325: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5326: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5327: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0080000000000:0:0:0:00:1:00800:
//------------------------

#2;
word <= 'h03f0080000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1333
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5328: ir 'h%h !== 'h0", ir); end	// Vector No: 1332
assert (op === 'h00) else begin fail = 1; $display("Error 5329: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5330: extop 'h%h !== 1", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 5331: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 03f0080000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0080000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1334
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5332: ir 'h%h !== 'h0", ir); end	// Vector No: 1333
assert (op === 'h00) else begin fail = 1; $display("Error 5333: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5334: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5335: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0080000000000:1:0:3:f0:0:00080:
//------------------------

#2;
word <= 'h03f0080000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1335
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5336: ir 'h%h !== 'h3", ir); end	// Vector No: 1334
assert (op === 'hf0) else begin fail = 1; $display("Error 5337: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5338: extop 'h%h !== 0", extop); end
assert (addr === 'h00080) else begin fail = 1; $display("Error 5339: addr 'h%h !== 'h00080", addr); end
#2;
clk <= 0;

// 03f0080000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0080000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1336
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5340: ir 'h%h !== 'h0", ir); end	// Vector No: 1335
assert (op === 'h00) else begin fail = 1; $display("Error 5341: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5342: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5343: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100003f00000:0:0:0:00:0:01000:
//------------------------

#2;
word <= 'h0000100003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1337
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5344: ir 'h%h !== 'h0", ir); end	// Vector No: 1336
assert (op === 'h00) else begin fail = 1; $display("Error 5345: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5346: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 5347: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 0000100003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000100003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1338
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5348: ir 'h%h !== 'h0", ir); end	// Vector No: 1337
assert (op === 'h00) else begin fail = 1; $display("Error 5349: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5350: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5351: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000100003f00000:1:0:0:00:0:00100:
//------------------------

#2;
word <= 'h0000100003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1339
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5352: ir 'h%h !== 'h0", ir); end	// Vector No: 1338
assert (op === 'h00) else begin fail = 1; $display("Error 5353: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5354: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 5355: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 0000100003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000100003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1340
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5356: ir 'h%h !== 'h0", ir); end	// Vector No: 1339
assert (op === 'h03) else begin fail = 1; $display("Error 5357: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5358: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5359: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0100000000000:0:0:0:01:1:01000:
//------------------------

#2;
word <= 'h03f0100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1341
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5360: ir 'h%h !== 'h0", ir); end	// Vector No: 1340
assert (op === 'h01) else begin fail = 1; $display("Error 5361: op 'h%h !== 'h01", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5362: extop 'h%h !== 1", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 5363: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 03f0100000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1342
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5364: ir 'h%h !== 'h0", ir); end	// Vector No: 1341
assert (op === 'h00) else begin fail = 1; $display("Error 5365: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5366: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5367: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0100000000000:1:0:3:f0:0:00100:
//------------------------

#2;
word <= 'h03f0100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1343
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5368: ir 'h%h !== 'h3", ir); end	// Vector No: 1342
assert (op === 'hf0) else begin fail = 1; $display("Error 5369: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5370: extop 'h%h !== 0", extop); end
assert (addr === 'h00100) else begin fail = 1; $display("Error 5371: addr 'h%h !== 'h00100", addr); end
#2;
clk <= 0;

// 03f0100000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1344
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5372: ir 'h%h !== 'h0", ir); end	// Vector No: 1343
assert (op === 'h00) else begin fail = 1; $display("Error 5373: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5374: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5375: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200003f00000:0:0:0:00:0:02000:
//------------------------

#2;
word <= 'h0000200003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1345
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5376: ir 'h%h !== 'h0", ir); end	// Vector No: 1344
assert (op === 'h00) else begin fail = 1; $display("Error 5377: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5378: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 5379: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 0000200003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000200003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1346
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5380: ir 'h%h !== 'h0", ir); end	// Vector No: 1345
assert (op === 'h00) else begin fail = 1; $display("Error 5381: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5382: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5383: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000200003f00000:1:0:0:00:0:00200:
//------------------------

#2;
word <= 'h0000200003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1347
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5384: ir 'h%h !== 'h0", ir); end	// Vector No: 1346
assert (op === 'h00) else begin fail = 1; $display("Error 5385: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5386: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 5387: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 0000200003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000200003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1348
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5388: ir 'h%h !== 'h0", ir); end	// Vector No: 1347
assert (op === 'h03) else begin fail = 1; $display("Error 5389: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5390: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5391: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0200000000000:0:0:0:02:1:02000:
//------------------------

#2;
word <= 'h03f0200000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1349
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5392: ir 'h%h !== 'h0", ir); end	// Vector No: 1348
assert (op === 'h02) else begin fail = 1; $display("Error 5393: op 'h%h !== 'h02", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5394: extop 'h%h !== 1", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 5395: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 03f0200000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0200000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1350
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5396: ir 'h%h !== 'h0", ir); end	// Vector No: 1349
assert (op === 'h00) else begin fail = 1; $display("Error 5397: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5398: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5399: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0200000000000:1:0:3:f0:0:00200:
//------------------------

#2;
word <= 'h03f0200000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1351
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5400: ir 'h%h !== 'h3", ir); end	// Vector No: 1350
assert (op === 'hf0) else begin fail = 1; $display("Error 5401: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5402: extop 'h%h !== 0", extop); end
assert (addr === 'h00200) else begin fail = 1; $display("Error 5403: addr 'h%h !== 'h00200", addr); end
#2;
clk <= 0;

// 03f0200000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0200000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1352
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5404: ir 'h%h !== 'h0", ir); end	// Vector No: 1351
assert (op === 'h00) else begin fail = 1; $display("Error 5405: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5406: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5407: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400003f00000:0:0:0:00:0:04000:
//------------------------

#2;
word <= 'h0000400003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1353
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5408: ir 'h%h !== 'h0", ir); end	// Vector No: 1352
assert (op === 'h00) else begin fail = 1; $display("Error 5409: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5410: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 5411: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 0000400003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000400003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1354
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5412: ir 'h%h !== 'h0", ir); end	// Vector No: 1353
assert (op === 'h00) else begin fail = 1; $display("Error 5413: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5414: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5415: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000400003f00000:1:0:0:00:0:00400:
//------------------------

#2;
word <= 'h0000400003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1355
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5416: ir 'h%h !== 'h0", ir); end	// Vector No: 1354
assert (op === 'h00) else begin fail = 1; $display("Error 5417: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5418: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 5419: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 0000400003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000400003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1356
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5420: ir 'h%h !== 'h0", ir); end	// Vector No: 1355
assert (op === 'h03) else begin fail = 1; $display("Error 5421: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5422: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5423: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0400000000000:0:0:0:04:1:04000:
//------------------------

#2;
word <= 'h03f0400000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1357
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5424: ir 'h%h !== 'h0", ir); end	// Vector No: 1356
assert (op === 'h04) else begin fail = 1; $display("Error 5425: op 'h%h !== 'h04", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5426: extop 'h%h !== 1", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 5427: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 03f0400000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0400000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1358
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5428: ir 'h%h !== 'h0", ir); end	// Vector No: 1357
assert (op === 'h00) else begin fail = 1; $display("Error 5429: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5430: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5431: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0400000000000:1:0:3:f0:0:00400:
//------------------------

#2;
word <= 'h03f0400000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1359
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5432: ir 'h%h !== 'h3", ir); end	// Vector No: 1358
assert (op === 'hf0) else begin fail = 1; $display("Error 5433: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5434: extop 'h%h !== 0", extop); end
assert (addr === 'h00400) else begin fail = 1; $display("Error 5435: addr 'h%h !== 'h00400", addr); end
#2;
clk <= 0;

// 03f0400000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0400000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1360
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5436: ir 'h%h !== 'h0", ir); end	// Vector No: 1359
assert (op === 'h00) else begin fail = 1; $display("Error 5437: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5438: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5439: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800003f00000:0:0:0:00:0:08000:
//------------------------

#2;
word <= 'h0000800003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1361
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5440: ir 'h%h !== 'h0", ir); end	// Vector No: 1360
assert (op === 'h00) else begin fail = 1; $display("Error 5441: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5442: extop 'h%h !== 0", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 5443: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 0000800003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0000800003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1362
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5444: ir 'h%h !== 'h0", ir); end	// Vector No: 1361
assert (op === 'h00) else begin fail = 1; $display("Error 5445: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5446: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5447: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0000800003f00000:1:0:0:00:0:00800:
//------------------------

#2;
word <= 'h0000800003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1363
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5448: ir 'h%h !== 'h0", ir); end	// Vector No: 1362
assert (op === 'h00) else begin fail = 1; $display("Error 5449: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5450: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 5451: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 0000800003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0000800003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1364
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5452: ir 'h%h !== 'h0", ir); end	// Vector No: 1363
assert (op === 'h03) else begin fail = 1; $display("Error 5453: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5454: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5455: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0800000000000:0:0:0:08:1:08000:
//------------------------

#2;
word <= 'h03f0800000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1365
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5456: ir 'h%h !== 'h0", ir); end	// Vector No: 1364
assert (op === 'h08) else begin fail = 1; $display("Error 5457: op 'h%h !== 'h08", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5458: extop 'h%h !== 1", extop); end
assert (addr === 'h08000) else begin fail = 1; $display("Error 5459: addr 'h%h !== 'h08000", addr); end
#2;
clk <= 0;

// 03f0800000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0800000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1366
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5460: ir 'h%h !== 'h0", ir); end	// Vector No: 1365
assert (op === 'h00) else begin fail = 1; $display("Error 5461: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5462: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5463: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0800000000000:1:0:3:f0:0:00800:
//------------------------

#2;
word <= 'h03f0800000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1367
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5464: ir 'h%h !== 'h3", ir); end	// Vector No: 1366
assert (op === 'hf0) else begin fail = 1; $display("Error 5465: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5466: extop 'h%h !== 0", extop); end
assert (addr === 'h00800) else begin fail = 1; $display("Error 5467: addr 'h%h !== 'h00800", addr); end
#2;
clk <= 0;

// 03f0800000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0800000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1368
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5468: ir 'h%h !== 'h0", ir); end	// Vector No: 1367
assert (op === 'h00) else begin fail = 1; $display("Error 5469: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5470: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5471: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000003f00000:0:0:0:00:0:10000:
//------------------------

#2;
word <= 'h0001000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1369
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5472: ir 'h%h !== 'h0", ir); end	// Vector No: 1368
assert (op === 'h00) else begin fail = 1; $display("Error 5473: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5474: extop 'h%h !== 0", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 5475: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 0001000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0001000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1370
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5476: ir 'h%h !== 'h0", ir); end	// Vector No: 1369
assert (op === 'h00) else begin fail = 1; $display("Error 5477: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5478: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5479: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000003f00000:1:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0001000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1371
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5480: ir 'h%h !== 'h0", ir); end	// Vector No: 1370
assert (op === 'h01) else begin fail = 1; $display("Error 5481: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5482: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5483: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0001000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0001000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1372
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5484: ir 'h%h !== 'h0", ir); end	// Vector No: 1371
assert (op === 'h03) else begin fail = 1; $display("Error 5485: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5486: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5487: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f1000000000000:0:0:0:10:1:10000:
//------------------------

#2;
word <= 'h03f1000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1373
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5488: ir 'h%h !== 'h0", ir); end	// Vector No: 1372
assert (op === 'h10) else begin fail = 1; $display("Error 5489: op 'h%h !== 'h10", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5490: extop 'h%h !== 1", extop); end
assert (addr === 'h10000) else begin fail = 1; $display("Error 5491: addr 'h%h !== 'h10000", addr); end
#2;
clk <= 0;

// 03f1000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f1000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1374
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5492: ir 'h%h !== 'h0", ir); end	// Vector No: 1373
assert (op === 'h00) else begin fail = 1; $display("Error 5493: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5494: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5495: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f1000000000000:1:0:3:f0:0:01000:
//------------------------

#2;
word <= 'h03f1000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1375
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5496: ir 'h%h !== 'h3", ir); end	// Vector No: 1374
assert (op === 'hf0) else begin fail = 1; $display("Error 5497: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5498: extop 'h%h !== 0", extop); end
assert (addr === 'h01000) else begin fail = 1; $display("Error 5499: addr 'h%h !== 'h01000", addr); end
#2;
clk <= 0;

// 03f1000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f1000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1376
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5500: ir 'h%h !== 'h0", ir); end	// Vector No: 1375
assert (op === 'h00) else begin fail = 1; $display("Error 5501: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5502: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5503: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000003f00000:0:0:0:00:0:20000:
//------------------------

#2;
word <= 'h0002000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1377
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5504: ir 'h%h !== 'h0", ir); end	// Vector No: 1376
assert (op === 'h00) else begin fail = 1; $display("Error 5505: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5506: extop 'h%h !== 0", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 5507: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 0002000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0002000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1378
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5508: ir 'h%h !== 'h0", ir); end	// Vector No: 1377
assert (op === 'h00) else begin fail = 1; $display("Error 5509: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5510: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5511: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000003f00000:1:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0002000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1379
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5512: ir 'h%h !== 'h0", ir); end	// Vector No: 1378
assert (op === 'h02) else begin fail = 1; $display("Error 5513: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5514: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5515: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0002000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0002000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1380
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5516: ir 'h%h !== 'h0", ir); end	// Vector No: 1379
assert (op === 'h03) else begin fail = 1; $display("Error 5517: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5518: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5519: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f2000000000000:0:0:0:20:1:20000:
//------------------------

#2;
word <= 'h03f2000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1381
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5520: ir 'h%h !== 'h0", ir); end	// Vector No: 1380
assert (op === 'h20) else begin fail = 1; $display("Error 5521: op 'h%h !== 'h20", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5522: extop 'h%h !== 1", extop); end
assert (addr === 'h20000) else begin fail = 1; $display("Error 5523: addr 'h%h !== 'h20000", addr); end
#2;
clk <= 0;

// 03f2000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f2000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1382
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5524: ir 'h%h !== 'h0", ir); end	// Vector No: 1381
assert (op === 'h00) else begin fail = 1; $display("Error 5525: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5526: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5527: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f2000000000000:1:0:3:f0:0:02000:
//------------------------

#2;
word <= 'h03f2000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1383
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5528: ir 'h%h !== 'h3", ir); end	// Vector No: 1382
assert (op === 'hf0) else begin fail = 1; $display("Error 5529: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5530: extop 'h%h !== 0", extop); end
assert (addr === 'h02000) else begin fail = 1; $display("Error 5531: addr 'h%h !== 'h02000", addr); end
#2;
clk <= 0;

// 03f2000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f2000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1384
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5532: ir 'h%h !== 'h0", ir); end	// Vector No: 1383
assert (op === 'h00) else begin fail = 1; $display("Error 5533: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5534: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5535: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000003f00000:0:0:0:00:0:40000:
//------------------------

#2;
word <= 'h0004000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1385
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5536: ir 'h%h !== 'h0", ir); end	// Vector No: 1384
assert (op === 'h00) else begin fail = 1; $display("Error 5537: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5538: extop 'h%h !== 0", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 5539: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 0004000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0004000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1386
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5540: ir 'h%h !== 'h0", ir); end	// Vector No: 1385
assert (op === 'h00) else begin fail = 1; $display("Error 5541: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5542: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5543: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000003f00000:1:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0004000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1387
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5544: ir 'h%h !== 'h0", ir); end	// Vector No: 1386
assert (op === 'h04) else begin fail = 1; $display("Error 5545: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5546: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5547: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0004000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0004000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1388
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5548: ir 'h%h !== 'h0", ir); end	// Vector No: 1387
assert (op === 'h03) else begin fail = 1; $display("Error 5549: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5550: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5551: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f4000000000000:0:0:0:40:1:40000:
//------------------------

#2;
word <= 'h03f4000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1389
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5552: ir 'h%h !== 'h0", ir); end	// Vector No: 1388
assert (op === 'h40) else begin fail = 1; $display("Error 5553: op 'h%h !== 'h40", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5554: extop 'h%h !== 1", extop); end
assert (addr === 'h40000) else begin fail = 1; $display("Error 5555: addr 'h%h !== 'h40000", addr); end
#2;
clk <= 0;

// 03f4000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f4000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1390
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5556: ir 'h%h !== 'h0", ir); end	// Vector No: 1389
assert (op === 'h00) else begin fail = 1; $display("Error 5557: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5558: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5559: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f4000000000000:1:0:3:f0:0:04000:
//------------------------

#2;
word <= 'h03f4000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1391
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5560: ir 'h%h !== 'h3", ir); end	// Vector No: 1390
assert (op === 'hf0) else begin fail = 1; $display("Error 5561: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5562: extop 'h%h !== 0", extop); end
assert (addr === 'h04000) else begin fail = 1; $display("Error 5563: addr 'h%h !== 'h04000", addr); end
#2;
clk <= 0;

// 03f4000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f4000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1392
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5564: ir 'h%h !== 'h0", ir); end	// Vector No: 1391
assert (op === 'h00) else begin fail = 1; $display("Error 5565: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5566: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5567: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000003f00000:0:0:0:00:0:80000:
//------------------------

#2;
word <= 'h0008000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1393
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5568: ir 'h%h !== 'h0", ir); end	// Vector No: 1392
assert (op === 'h00) else begin fail = 1; $display("Error 5569: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5570: extop 'h%h !== 0", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 5571: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 0008000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0008000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1394
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5572: ir 'h%h !== 'h0", ir); end	// Vector No: 1393
assert (op === 'h00) else begin fail = 1; $display("Error 5573: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5574: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5575: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000003f00000:1:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0008000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1395
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5576: ir 'h%h !== 'h0", ir); end	// Vector No: 1394
assert (op === 'h08) else begin fail = 1; $display("Error 5577: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5578: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5579: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0008000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0008000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1396
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5580: ir 'h%h !== 'h0", ir); end	// Vector No: 1395
assert (op === 'h03) else begin fail = 1; $display("Error 5581: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5582: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5583: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f8000000000000:0:0:0:80:1:80000:
//------------------------

#2;
word <= 'h03f8000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1397
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5584: ir 'h%h !== 'h0", ir); end	// Vector No: 1396
assert (op === 'h80) else begin fail = 1; $display("Error 5585: op 'h%h !== 'h80", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5586: extop 'h%h !== 1", extop); end
assert (addr === 'h80000) else begin fail = 1; $display("Error 5587: addr 'h%h !== 'h80000", addr); end
#2;
clk <= 0;

// 03f8000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f8000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1398
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5588: ir 'h%h !== 'h0", ir); end	// Vector No: 1397
assert (op === 'h00) else begin fail = 1; $display("Error 5589: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5590: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5591: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f8000000000000:1:0:3:f8:0:00000:
//------------------------

#2;
word <= 'h03f8000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1399
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5592: ir 'h%h !== 'h3", ir); end	// Vector No: 1398
assert (op === 'hf8) else begin fail = 1; $display("Error 5593: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5594: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5595: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f8000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f8000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1400
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5596: ir 'h%h !== 'h0", ir); end	// Vector No: 1399
assert (op === 'h00) else begin fail = 1; $display("Error 5597: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5598: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5599: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000003f00000:0:0:0:01:0:00000:
//------------------------

#2;
word <= 'h0010000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1401
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5600: ir 'h%h !== 'h0", ir); end	// Vector No: 1400
assert (op === 'h01) else begin fail = 1; $display("Error 5601: op 'h%h !== 'h01", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5602: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5603: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0010000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1402
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5604: ir 'h%h !== 'h0", ir); end	// Vector No: 1401
assert (op === 'h00) else begin fail = 1; $display("Error 5605: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5606: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5607: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000003f00000:1:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0010000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1403
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5608: ir 'h%h !== 'h0", ir); end	// Vector No: 1402
assert (op === 'h10) else begin fail = 1; $display("Error 5609: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5610: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5611: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0010000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0010000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1404
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5612: ir 'h%h !== 'h0", ir); end	// Vector No: 1403
assert (op === 'h03) else begin fail = 1; $display("Error 5613: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5614: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5615: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 03f0000000000000:0:0:0:00:1:00000:
//------------------------

#2;
word <= 'h03f0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1405
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5616: ir 'h%h !== 'h0", ir); end	// Vector No: 1404
assert (op === 'h00) else begin fail = 1; $display("Error 5617: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5618: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5619: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1406
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5620: ir 'h%h !== 'h0", ir); end	// Vector No: 1405
assert (op === 'h00) else begin fail = 1; $display("Error 5621: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5622: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5623: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h03f0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1407
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5624: ir 'h%h !== 'h3", ir); end	// Vector No: 1406
assert (op === 'hf0) else begin fail = 1; $display("Error 5625: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5626: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5627: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 03f0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h03f0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1408
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5628: ir 'h%h !== 'h0", ir); end	// Vector No: 1407
assert (op === 'h00) else begin fail = 1; $display("Error 5629: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5630: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5631: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000003f00000:0:0:0:02:0:00000:
//------------------------

#2;
word <= 'h0020000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1409
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5632: ir 'h%h !== 'h0", ir); end	// Vector No: 1408
assert (op === 'h02) else begin fail = 1; $display("Error 5633: op 'h%h !== 'h02", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5634: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5635: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0020000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1410
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5636: ir 'h%h !== 'h0", ir); end	// Vector No: 1409
assert (op === 'h00) else begin fail = 1; $display("Error 5637: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5638: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5639: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000003f00000:1:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0020000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1411
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5640: ir 'h%h !== 'h0", ir); end	// Vector No: 1410
assert (op === 'h20) else begin fail = 1; $display("Error 5641: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5642: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5643: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0020000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0020000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1412
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5644: ir 'h%h !== 'h0", ir); end	// Vector No: 1411
assert (op === 'h03) else begin fail = 1; $display("Error 5645: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5646: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5647: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0040000003f00000:0:0:0:04:0:00000:
//------------------------

#2;
word <= 'h0040000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1413
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5648: ir 'h%h !== 'h0", ir); end	// Vector No: 1412
assert (op === 'h04) else begin fail = 1; $display("Error 5649: op 'h%h !== 'h04", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5650: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5651: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0040000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1414
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5652: ir 'h%h !== 'h0", ir); end	// Vector No: 1413
assert (op === 'h00) else begin fail = 1; $display("Error 5653: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5654: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5655: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0040000003f00000:1:0:0:40:0:07000:
//------------------------

#2;
word <= 'h0040000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1415
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5656: ir 'h%h !== 'h0", ir); end	// Vector No: 1414
assert (op === 'h40) else begin fail = 1; $display("Error 5657: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5658: extop 'h%h !== 0", extop); end
assert (addr === 'h07000) else begin fail = 1; $display("Error 5659: addr 'h%h !== 'h07000", addr); end
#2;
clk <= 0;

// 0040000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0040000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1416
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5660: ir 'h%h !== 'h0", ir); end	// Vector No: 1415
assert (op === 'h03) else begin fail = 1; $display("Error 5661: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5662: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5663: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0080000003f00000:0:0:0:08:0:00000:
//------------------------

#2;
word <= 'h0080000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1417
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5664: ir 'h%h !== 'h0", ir); end	// Vector No: 1416
assert (op === 'h08) else begin fail = 1; $display("Error 5665: op 'h%h !== 'h08", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5666: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5667: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0080000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1418
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5668: ir 'h%h !== 'h0", ir); end	// Vector No: 1417
assert (op === 'h00) else begin fail = 1; $display("Error 5669: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5670: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5671: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000003f00000:1:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0080000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1419
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5672: ir 'h%h !== 'h0", ir); end	// Vector No: 1418
assert (op === 'h80) else begin fail = 1; $display("Error 5673: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5674: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5675: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0080000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0080000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1420
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5676: ir 'h%h !== 'h0", ir); end	// Vector No: 1419
assert (op === 'h03) else begin fail = 1; $display("Error 5677: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5678: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5679: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0100000003f00000:0:0:0:10:0:00000:
//------------------------

#2;
word <= 'h0100000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1421
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5680: ir 'h%h !== 'h0", ir); end	// Vector No: 1420
assert (op === 'h10) else begin fail = 1; $display("Error 5681: op 'h%h !== 'h10", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5682: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5683: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0100000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1422
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5684: ir 'h%h !== 'h0", ir); end	// Vector No: 1421
assert (op === 'h00) else begin fail = 1; $display("Error 5685: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5686: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5687: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000003f00000:1:0:1:00:0:00000:
//------------------------

#2;
word <= 'h0100000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1423
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 5688: ir 'h%h !== 'h1", ir); end	// Vector No: 1422
assert (op === 'h00) else begin fail = 1; $display("Error 5689: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5690: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5691: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0100000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0100000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1424
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5692: ir 'h%h !== 'h0", ir); end	// Vector No: 1423
assert (op === 'h03) else begin fail = 1; $display("Error 5693: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5694: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5695: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0200000003f00000:0:0:0:20:0:00000:
//------------------------

#2;
word <= 'h0200000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1425
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5696: ir 'h%h !== 'h0", ir); end	// Vector No: 1424
assert (op === 'h20) else begin fail = 1; $display("Error 5697: op 'h%h !== 'h20", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5698: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5699: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0200000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1426
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5700: ir 'h%h !== 'h0", ir); end	// Vector No: 1425
assert (op === 'h00) else begin fail = 1; $display("Error 5701: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5702: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5703: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000003f00000:1:0:2:00:0:00000:
//------------------------

#2;
word <= 'h0200000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1427
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 5704: ir 'h%h !== 'h2", ir); end	// Vector No: 1426
assert (op === 'h00) else begin fail = 1; $display("Error 5705: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5706: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5707: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0200000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0200000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1428
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5708: ir 'h%h !== 'h0", ir); end	// Vector No: 1427
assert (op === 'h03) else begin fail = 1; $display("Error 5709: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5710: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5711: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0400000003f00000:0:0:0:40:0:00000:
//------------------------

#2;
word <= 'h0400000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1429
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5712: ir 'h%h !== 'h0", ir); end	// Vector No: 1428
assert (op === 'h40) else begin fail = 1; $display("Error 5713: op 'h%h !== 'h40", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5714: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5715: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0400000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1430
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5716: ir 'h%h !== 'h0", ir); end	// Vector No: 1429
assert (op === 'h00) else begin fail = 1; $display("Error 5717: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5718: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5719: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000003f00000:1:0:4:00:0:00000:
//------------------------

#2;
word <= 'h0400000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1431
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 5720: ir 'h%h !== 'h4", ir); end	// Vector No: 1430
assert (op === 'h00) else begin fail = 1; $display("Error 5721: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5722: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5723: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0400000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0400000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1432
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5724: ir 'h%h !== 'h0", ir); end	// Vector No: 1431
assert (op === 'h03) else begin fail = 1; $display("Error 5725: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5726: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5727: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 0800000003f00000:0:0:0:80:0:00000:
//------------------------

#2;
word <= 'h0800000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1433
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5728: ir 'h%h !== 'h0", ir); end	// Vector No: 1432
assert (op === 'h80) else begin fail = 1; $display("Error 5729: op 'h%h !== 'h80", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5730: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5731: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h0800000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1434
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5732: ir 'h%h !== 'h0", ir); end	// Vector No: 1433
assert (op === 'h00) else begin fail = 1; $display("Error 5733: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5734: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5735: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000003f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h0800000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1435
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5736: ir 'h%h !== 'h0", ir); end	// Vector No: 1434
assert (op === 'h00) else begin fail = 1; $display("Error 5737: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5738: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5739: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 0800000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h0800000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1436
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5740: ir 'h%h !== 'h0", ir); end	// Vector No: 1435
assert (op === 'h03) else begin fail = 1; $display("Error 5741: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5742: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5743: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 1000000003f00000:0:0:1:00:0:00000:
//------------------------

#2;
word <= 'h1000000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1437
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 5744: ir 'h%h !== 'h1", ir); end	// Vector No: 1436
assert (op === 'h00) else begin fail = 1; $display("Error 5745: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5746: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5747: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h1000000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1438
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5748: ir 'h%h !== 'h0", ir); end	// Vector No: 1437
assert (op === 'h00) else begin fail = 1; $display("Error 5749: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5750: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5751: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000003f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h1000000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1439
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5752: ir 'h%h !== 'h0", ir); end	// Vector No: 1438
assert (op === 'h00) else begin fail = 1; $display("Error 5753: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5754: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5755: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 1000000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h1000000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1440
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5756: ir 'h%h !== 'h0", ir); end	// Vector No: 1439
assert (op === 'h03) else begin fail = 1; $display("Error 5757: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5758: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5759: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 13f0000000000000:0:0:1:00:1:00000:
//------------------------

#2;
word <= 'h13f0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1441
#2;

assert (ir === 'h1) else begin fail = 1; $display("Error 5760: ir 'h%h !== 'h1", ir); end	// Vector No: 1440
assert (op === 'h00) else begin fail = 1; $display("Error 5761: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5762: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5763: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 13f0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h13f0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1442
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5764: ir 'h%h !== 'h0", ir); end	// Vector No: 1441
assert (op === 'h00) else begin fail = 1; $display("Error 5765: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5766: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5767: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 13f0000000000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h13f0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1443
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5768: ir 'h%h !== 'h3", ir); end	// Vector No: 1442
assert (op === 'hf0) else begin fail = 1; $display("Error 5769: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5770: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5771: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 13f0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h13f0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1444
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5772: ir 'h%h !== 'h0", ir); end	// Vector No: 1443
assert (op === 'h00) else begin fail = 1; $display("Error 5773: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5774: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5775: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000003f00000:0:0:2:00:0:00000:
//------------------------

#2;
word <= 'h2000000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1445
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 5776: ir 'h%h !== 'h2", ir); end	// Vector No: 1444
assert (op === 'h00) else begin fail = 1; $display("Error 5777: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5778: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5779: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h2000000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1446
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5780: ir 'h%h !== 'h0", ir); end	// Vector No: 1445
assert (op === 'h00) else begin fail = 1; $display("Error 5781: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5782: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5783: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000003f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h2000000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1447
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5784: ir 'h%h !== 'h0", ir); end	// Vector No: 1446
assert (op === 'h00) else begin fail = 1; $display("Error 5785: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5786: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5787: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 2000000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h2000000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1448
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5788: ir 'h%h !== 'h0", ir); end	// Vector No: 1447
assert (op === 'h03) else begin fail = 1; $display("Error 5789: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5790: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5791: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 23f0000000000000:0:0:2:00:1:00000:
//------------------------

#2;
word <= 'h23f0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1449
#2;

assert (ir === 'h2) else begin fail = 1; $display("Error 5792: ir 'h%h !== 'h2", ir); end	// Vector No: 1448
assert (op === 'h00) else begin fail = 1; $display("Error 5793: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5794: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5795: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 23f0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h23f0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1450
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5796: ir 'h%h !== 'h0", ir); end	// Vector No: 1449
assert (op === 'h00) else begin fail = 1; $display("Error 5797: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5798: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5799: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 23f0000000000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h23f0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1451
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5800: ir 'h%h !== 'h3", ir); end	// Vector No: 1450
assert (op === 'hf0) else begin fail = 1; $display("Error 5801: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5802: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5803: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 23f0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h23f0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1452
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5804: ir 'h%h !== 'h0", ir); end	// Vector No: 1451
assert (op === 'h00) else begin fail = 1; $display("Error 5805: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5806: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5807: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000003f00000:0:0:4:00:0:00000:
//------------------------

#2;
word <= 'h4000000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1453
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 5808: ir 'h%h !== 'h4", ir); end	// Vector No: 1452
assert (op === 'h00) else begin fail = 1; $display("Error 5809: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5810: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5811: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h4000000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1454
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5812: ir 'h%h !== 'h0", ir); end	// Vector No: 1453
assert (op === 'h00) else begin fail = 1; $display("Error 5813: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5814: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5815: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000003f00000:1:0:0:00:0:00000:
//------------------------

#2;
word <= 'h4000000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1455
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5816: ir 'h%h !== 'h0", ir); end	// Vector No: 1454
assert (op === 'h00) else begin fail = 1; $display("Error 5817: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5818: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5819: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 4000000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h4000000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1456
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5820: ir 'h%h !== 'h0", ir); end	// Vector No: 1455
assert (op === 'h03) else begin fail = 1; $display("Error 5821: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5822: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5823: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 43f0000000000000:0:0:4:00:1:00000:
//------------------------

#2;
word <= 'h43f0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1457
#2;

assert (ir === 'h4) else begin fail = 1; $display("Error 5824: ir 'h%h !== 'h4", ir); end	// Vector No: 1456
assert (op === 'h00) else begin fail = 1; $display("Error 5825: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5826: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5827: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 43f0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h43f0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1458
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5828: ir 'h%h !== 'h0", ir); end	// Vector No: 1457
assert (op === 'h00) else begin fail = 1; $display("Error 5829: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5830: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5831: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 43f0000000000000:1:0:3:f0:0:00000:
//------------------------

#2;
word <= 'h43f0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1459
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 5832: ir 'h%h !== 'h3", ir); end	// Vector No: 1458
assert (op === 'hf0) else begin fail = 1; $display("Error 5833: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5834: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5835: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 43f0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h43f0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1460
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5836: ir 'h%h !== 'h0", ir); end	// Vector No: 1459
assert (op === 'h00) else begin fail = 1; $display("Error 5837: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5838: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5839: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000003f00000:0:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000003f00000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1461
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 5840: ir 'h%h !== 'h8", ir); end	// Vector No: 1460
assert (op === 'h00) else begin fail = 1; $display("Error 5841: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5842: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5843: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000003f00000:0:1:0:00:1:00000:
//------------------------

#2;
word <= 'h8000000003f00000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1462
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5844: ir 'h%h !== 'h0", ir); end	// Vector No: 1461
assert (op === 'h00) else begin fail = 1; $display("Error 5845: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5846: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5847: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000003f00000:1:0:8:00:0:00000:
//------------------------

#2;
word <= 'h8000000003f00000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1463
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 5848: ir 'h%h !== 'h8", ir); end	// Vector No: 1462
assert (op === 'h00) else begin fail = 1; $display("Error 5849: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5850: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5851: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 8000000003f00000:1:1:0:03:0:00f00:
//------------------------

#2;
word <= 'h8000000003f00000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1464
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5852: ir 'h%h !== 'h0", ir); end	// Vector No: 1463
assert (op === 'h03) else begin fail = 1; $display("Error 5853: op 'h%h !== 'h03", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5854: extop 'h%h !== 0", extop); end
assert (addr === 'h00f00) else begin fail = 1; $display("Error 5855: addr 'h%h !== 'h00f00", addr); end
#2;
clk <= 0;

// 83f0000000000000:0:0:8:00:1:00000:
//------------------------

#2;
word <= 'h83f0000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1465
#2;

assert (ir === 'h8) else begin fail = 1; $display("Error 5856: ir 'h%h !== 'h8", ir); end	// Vector No: 1464
assert (op === 'h00) else begin fail = 1; $display("Error 5857: op 'h%h !== 'h00", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5858: extop 'h%h !== 1", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5859: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 83f0000000000000:0:1:0:00:0:00000:
//------------------------

#2;
word <= 'h83f0000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1466
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5860: ir 'h%h !== 'h0", ir); end	// Vector No: 1465
assert (op === 'h00) else begin fail = 1; $display("Error 5861: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5862: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5863: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 83f0000000000000:1:0:b:f0:0:00000:
//------------------------

#2;
word <= 'h83f0000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1467
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 5864: ir 'h%h !== 'hb", ir); end	// Vector No: 1466
assert (op === 'hf0) else begin fail = 1; $display("Error 5865: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5866: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5867: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// 83f0000000000000:1:1:0:00:0:00000:
//------------------------

#2;
word <= 'h83f0000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1468
#2;

assert (ir === 'h0) else begin fail = 1; $display("Error 5868: ir 'h%h !== 'h0", ir); end	// Vector No: 1467
assert (op === 'h00) else begin fail = 1; $display("Error 5869: op 'h%h !== 'h00", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5870: extop 'h%h !== 0", extop); end
assert (addr === 'h00000) else begin fail = 1; $display("Error 5871: addr 'h%h !== 'h00000", addr); end
#2;
clk <= 0;

// fffffffff3fffffe:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffffe;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1469
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5872: ir 'h%h !== 'hf", ir); end	// Vector No: 1468
assert (op === 'hff) else begin fail = 1; $display("Error 5873: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5874: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5875: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffffe:0:1:f:ff:1:ffffe:
//------------------------

#2;
word <= 'hfffffffff3fffffe;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1470
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5876: ir 'h%h !== 'hf", ir); end	// Vector No: 1469
assert (op === 'hff) else begin fail = 1; $display("Error 5877: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5878: extop 'h%h !== 1", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 5879: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// fffffffff3fffffe:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffffe;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1471
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5880: ir 'h%h !== 'hf", ir); end	// Vector No: 1470
assert (op === 'hf8) else begin fail = 1; $display("Error 5881: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5882: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5883: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffffe:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffffe;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1472
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5884: ir 'h%h !== 'hf", ir); end	// Vector No: 1471
assert (op === 'hf0) else begin fail = 1; $display("Error 5885: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5886: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 5887: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffe:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffffe;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1473
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5888: ir 'h%h !== 'hf", ir); end	// Vector No: 1472
assert (op === 'hff) else begin fail = 1; $display("Error 5889: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5890: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5891: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffffe:0:1:f:ff:0:ffffe:
//------------------------

#2;
word <= 'hf3fffffffffffffe;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1474
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5892: ir 'h%h !== 'hf", ir); end	// Vector No: 1473
assert (op === 'hff) else begin fail = 1; $display("Error 5893: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5894: extop 'h%h !== 0", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 5895: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// f3fffffffffffffe:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffe;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1475
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 5896: ir 'h%h !== 'hb", ir); end	// Vector No: 1474
assert (op === 'hf8) else begin fail = 1; $display("Error 5897: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5898: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5899: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffe:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffe;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1476
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5900: ir 'h%h !== 'hf", ir); end	// Vector No: 1475
assert (op === 'hf8) else begin fail = 1; $display("Error 5901: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5902: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5903: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffffd:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffffd;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1477
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5904: ir 'h%h !== 'hf", ir); end	// Vector No: 1476
assert (op === 'hff) else begin fail = 1; $display("Error 5905: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5906: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5907: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffffd:0:1:f:ff:1:ffffd:
//------------------------

#2;
word <= 'hfffffffff3fffffd;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1478
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5908: ir 'h%h !== 'hf", ir); end	// Vector No: 1477
assert (op === 'hff) else begin fail = 1; $display("Error 5909: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5910: extop 'h%h !== 1", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 5911: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// fffffffff3fffffd:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffffd;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1479
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5912: ir 'h%h !== 'hf", ir); end	// Vector No: 1478
assert (op === 'hf8) else begin fail = 1; $display("Error 5913: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5914: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5915: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffffd:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffffd;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1480
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5916: ir 'h%h !== 'hf", ir); end	// Vector No: 1479
assert (op === 'hf0) else begin fail = 1; $display("Error 5917: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5918: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 5919: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffd:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffffd;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1481
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5920: ir 'h%h !== 'hf", ir); end	// Vector No: 1480
assert (op === 'hff) else begin fail = 1; $display("Error 5921: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5922: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5923: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffffd:0:1:f:ff:0:ffffd:
//------------------------

#2;
word <= 'hf3fffffffffffffd;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1482
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5924: ir 'h%h !== 'hf", ir); end	// Vector No: 1481
assert (op === 'hff) else begin fail = 1; $display("Error 5925: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5926: extop 'h%h !== 0", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 5927: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// f3fffffffffffffd:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffd;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1483
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 5928: ir 'h%h !== 'hb", ir); end	// Vector No: 1482
assert (op === 'hf8) else begin fail = 1; $display("Error 5929: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5930: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5931: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffd:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffd;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1484
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5932: ir 'h%h !== 'hf", ir); end	// Vector No: 1483
assert (op === 'hf8) else begin fail = 1; $display("Error 5933: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5934: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5935: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffffb:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffffb;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1485
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5936: ir 'h%h !== 'hf", ir); end	// Vector No: 1484
assert (op === 'hff) else begin fail = 1; $display("Error 5937: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5938: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5939: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffffb:0:1:f:ff:1:ffffb:
//------------------------

#2;
word <= 'hfffffffff3fffffb;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1486
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5940: ir 'h%h !== 'hf", ir); end	// Vector No: 1485
assert (op === 'hff) else begin fail = 1; $display("Error 5941: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5942: extop 'h%h !== 1", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 5943: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// fffffffff3fffffb:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffffb;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1487
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5944: ir 'h%h !== 'hf", ir); end	// Vector No: 1486
assert (op === 'hf8) else begin fail = 1; $display("Error 5945: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5946: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5947: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffffb:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffffb;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1488
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5948: ir 'h%h !== 'hf", ir); end	// Vector No: 1487
assert (op === 'hf0) else begin fail = 1; $display("Error 5949: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5950: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 5951: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffb:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffffb;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1489
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5952: ir 'h%h !== 'hf", ir); end	// Vector No: 1488
assert (op === 'hff) else begin fail = 1; $display("Error 5953: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5954: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5955: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffffb:0:1:f:ff:0:ffffb:
//------------------------

#2;
word <= 'hf3fffffffffffffb;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1490
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5956: ir 'h%h !== 'hf", ir); end	// Vector No: 1489
assert (op === 'hff) else begin fail = 1; $display("Error 5957: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5958: extop 'h%h !== 0", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 5959: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// f3fffffffffffffb:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffb;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1491
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 5960: ir 'h%h !== 'hb", ir); end	// Vector No: 1490
assert (op === 'hf8) else begin fail = 1; $display("Error 5961: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5962: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5963: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffffb:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffffb;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1492
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5964: ir 'h%h !== 'hf", ir); end	// Vector No: 1491
assert (op === 'hf8) else begin fail = 1; $display("Error 5965: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5966: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5967: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffff7:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffff7;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1493
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5968: ir 'h%h !== 'hf", ir); end	// Vector No: 1492
assert (op === 'hff) else begin fail = 1; $display("Error 5969: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5970: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5971: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffff7:0:1:f:ff:1:ffff7:
//------------------------

#2;
word <= 'hfffffffff3fffff7;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1494
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5972: ir 'h%h !== 'hf", ir); end	// Vector No: 1493
assert (op === 'hff) else begin fail = 1; $display("Error 5973: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5974: extop 'h%h !== 1", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 5975: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// fffffffff3fffff7:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffff7;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1495
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5976: ir 'h%h !== 'hf", ir); end	// Vector No: 1494
assert (op === 'hf8) else begin fail = 1; $display("Error 5977: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5978: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5979: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffff7:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffff7;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1496
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5980: ir 'h%h !== 'hf", ir); end	// Vector No: 1495
assert (op === 'hf0) else begin fail = 1; $display("Error 5981: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5982: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 5983: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffff7:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffff7;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1497
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5984: ir 'h%h !== 'hf", ir); end	// Vector No: 1496
assert (op === 'hff) else begin fail = 1; $display("Error 5985: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 5986: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 5987: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffff7:0:1:f:ff:0:ffff7:
//------------------------

#2;
word <= 'hf3fffffffffffff7;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1498
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5988: ir 'h%h !== 'hf", ir); end	// Vector No: 1497
assert (op === 'hff) else begin fail = 1; $display("Error 5989: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5990: extop 'h%h !== 0", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 5991: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// f3fffffffffffff7:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffff7;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1499
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 5992: ir 'h%h !== 'hb", ir); end	// Vector No: 1498
assert (op === 'hf8) else begin fail = 1; $display("Error 5993: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5994: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5995: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffff7:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffff7;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1500
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 5996: ir 'h%h !== 'hf", ir); end	// Vector No: 1499
assert (op === 'hf8) else begin fail = 1; $display("Error 5997: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 5998: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 5999: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffef:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffffef;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1501
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6000: ir 'h%h !== 'hf", ir); end	// Vector No: 1500
assert (op === 'hff) else begin fail = 1; $display("Error 6001: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6002: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6003: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffffef:0:1:f:ff:1:fffef:
//------------------------

#2;
word <= 'hfffffffff3ffffef;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1502
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6004: ir 'h%h !== 'hf", ir); end	// Vector No: 1501
assert (op === 'hff) else begin fail = 1; $display("Error 6005: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6006: extop 'h%h !== 1", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 6007: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// fffffffff3ffffef:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffffef;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1503
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6008: ir 'h%h !== 'hf", ir); end	// Vector No: 1502
assert (op === 'hf8) else begin fail = 1; $display("Error 6009: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6010: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6011: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffef:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3ffffef;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1504
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6012: ir 'h%h !== 'hf", ir); end	// Vector No: 1503
assert (op === 'hf0) else begin fail = 1; $display("Error 6013: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6014: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6015: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffef:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffffef;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1505
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6016: ir 'h%h !== 'hf", ir); end	// Vector No: 1504
assert (op === 'hff) else begin fail = 1; $display("Error 6017: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6018: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6019: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffffef:0:1:f:ff:0:fffef:
//------------------------

#2;
word <= 'hf3ffffffffffffef;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1506
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6020: ir 'h%h !== 'hf", ir); end	// Vector No: 1505
assert (op === 'hff) else begin fail = 1; $display("Error 6021: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6022: extop 'h%h !== 0", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 6023: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// f3ffffffffffffef:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffef;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1507
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6024: ir 'h%h !== 'hb", ir); end	// Vector No: 1506
assert (op === 'hf8) else begin fail = 1; $display("Error 6025: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6026: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6027: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffef:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffef;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1508
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6028: ir 'h%h !== 'hf", ir); end	// Vector No: 1507
assert (op === 'hf8) else begin fail = 1; $display("Error 6029: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6030: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6031: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffdf:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffffdf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1509
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6032: ir 'h%h !== 'hf", ir); end	// Vector No: 1508
assert (op === 'hff) else begin fail = 1; $display("Error 6033: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6034: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6035: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffffdf:0:1:f:ff:1:fffdf:
//------------------------

#2;
word <= 'hfffffffff3ffffdf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1510
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6036: ir 'h%h !== 'hf", ir); end	// Vector No: 1509
assert (op === 'hff) else begin fail = 1; $display("Error 6037: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6038: extop 'h%h !== 1", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 6039: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// fffffffff3ffffdf:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffffdf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1511
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6040: ir 'h%h !== 'hf", ir); end	// Vector No: 1510
assert (op === 'hf8) else begin fail = 1; $display("Error 6041: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6042: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6043: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffdf:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3ffffdf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1512
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6044: ir 'h%h !== 'hf", ir); end	// Vector No: 1511
assert (op === 'hf0) else begin fail = 1; $display("Error 6045: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6046: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6047: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffdf:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffffdf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1513
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6048: ir 'h%h !== 'hf", ir); end	// Vector No: 1512
assert (op === 'hff) else begin fail = 1; $display("Error 6049: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6050: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6051: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffffdf:0:1:f:ff:0:fffdf:
//------------------------

#2;
word <= 'hf3ffffffffffffdf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1514
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6052: ir 'h%h !== 'hf", ir); end	// Vector No: 1513
assert (op === 'hff) else begin fail = 1; $display("Error 6053: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6054: extop 'h%h !== 0", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 6055: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// f3ffffffffffffdf:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffdf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1515
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6056: ir 'h%h !== 'hb", ir); end	// Vector No: 1514
assert (op === 'hf8) else begin fail = 1; $display("Error 6057: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6058: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6059: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffdf:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffdf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1516
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6060: ir 'h%h !== 'hf", ir); end	// Vector No: 1515
assert (op === 'hf8) else begin fail = 1; $display("Error 6061: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6062: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6063: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffbf:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffffbf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1517
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6064: ir 'h%h !== 'hf", ir); end	// Vector No: 1516
assert (op === 'hff) else begin fail = 1; $display("Error 6065: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6066: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6067: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffffbf:0:1:f:ff:1:fffbf:
//------------------------

#2;
word <= 'hfffffffff3ffffbf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1518
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6068: ir 'h%h !== 'hf", ir); end	// Vector No: 1517
assert (op === 'hff) else begin fail = 1; $display("Error 6069: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6070: extop 'h%h !== 1", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 6071: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// fffffffff3ffffbf:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffffbf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1519
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6072: ir 'h%h !== 'hf", ir); end	// Vector No: 1518
assert (op === 'hf8) else begin fail = 1; $display("Error 6073: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6074: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6075: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffbf:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3ffffbf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1520
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6076: ir 'h%h !== 'hf", ir); end	// Vector No: 1519
assert (op === 'hf0) else begin fail = 1; $display("Error 6077: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6078: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6079: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffbf:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffffbf;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1521
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6080: ir 'h%h !== 'hf", ir); end	// Vector No: 1520
assert (op === 'hff) else begin fail = 1; $display("Error 6081: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6082: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6083: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffffbf:0:1:f:ff:0:fffbf:
//------------------------

#2;
word <= 'hf3ffffffffffffbf;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1522
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6084: ir 'h%h !== 'hf", ir); end	// Vector No: 1521
assert (op === 'hff) else begin fail = 1; $display("Error 6085: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6086: extop 'h%h !== 0", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 6087: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// f3ffffffffffffbf:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffbf;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1523
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6088: ir 'h%h !== 'hb", ir); end	// Vector No: 1522
assert (op === 'hf8) else begin fail = 1; $display("Error 6089: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6090: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6091: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffbf:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffbf;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1524
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6092: ir 'h%h !== 'hf", ir); end	// Vector No: 1523
assert (op === 'hf8) else begin fail = 1; $display("Error 6093: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6094: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6095: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffff7f:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffff7f;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1525
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6096: ir 'h%h !== 'hf", ir); end	// Vector No: 1524
assert (op === 'hff) else begin fail = 1; $display("Error 6097: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6098: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6099: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffff7f:0:1:f:ff:1:fff7f:
//------------------------

#2;
word <= 'hfffffffff3ffff7f;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1526
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6100: ir 'h%h !== 'hf", ir); end	// Vector No: 1525
assert (op === 'hff) else begin fail = 1; $display("Error 6101: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6102: extop 'h%h !== 1", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 6103: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// fffffffff3ffff7f:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffff7f;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1527
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6104: ir 'h%h !== 'hf", ir); end	// Vector No: 1526
assert (op === 'hf8) else begin fail = 1; $display("Error 6105: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6106: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6107: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffff7f:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3ffff7f;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1528
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6108: ir 'h%h !== 'hf", ir); end	// Vector No: 1527
assert (op === 'hf0) else begin fail = 1; $display("Error 6109: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6110: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6111: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffffff7f:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffff7f;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1529
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6112: ir 'h%h !== 'hf", ir); end	// Vector No: 1528
assert (op === 'hff) else begin fail = 1; $display("Error 6113: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6114: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6115: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffff7f:0:1:f:ff:0:fff7f:
//------------------------

#2;
word <= 'hf3ffffffffffff7f;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1530
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6116: ir 'h%h !== 'hf", ir); end	// Vector No: 1529
assert (op === 'hff) else begin fail = 1; $display("Error 6117: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6118: extop 'h%h !== 0", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 6119: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// f3ffffffffffff7f:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffff7f;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1531
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6120: ir 'h%h !== 'hb", ir); end	// Vector No: 1530
assert (op === 'hf8) else begin fail = 1; $display("Error 6121: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6122: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6123: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffff7f:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffff7f;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1532
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6124: ir 'h%h !== 'hf", ir); end	// Vector No: 1531
assert (op === 'hf8) else begin fail = 1; $display("Error 6125: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6126: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6127: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffeff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffeff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1533
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6128: ir 'h%h !== 'hf", ir); end	// Vector No: 1532
assert (op === 'hff) else begin fail = 1; $display("Error 6129: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6130: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6131: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffeff:0:1:f:ff:1:ffeff:
//------------------------

#2;
word <= 'hfffffffff3fffeff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1534
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6132: ir 'h%h !== 'hf", ir); end	// Vector No: 1533
assert (op === 'hff) else begin fail = 1; $display("Error 6133: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6134: extop 'h%h !== 1", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 6135: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// fffffffff3fffeff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffeff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1535
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6136: ir 'h%h !== 'hf", ir); end	// Vector No: 1534
assert (op === 'hf8) else begin fail = 1; $display("Error 6137: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6138: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6139: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffeff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffeff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1536
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6140: ir 'h%h !== 'hf", ir); end	// Vector No: 1535
assert (op === 'hf0) else begin fail = 1; $display("Error 6141: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6142: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6143: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffeff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffeff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1537
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6144: ir 'h%h !== 'hf", ir); end	// Vector No: 1536
assert (op === 'hff) else begin fail = 1; $display("Error 6145: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6146: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6147: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffeff:0:1:f:ff:0:ffeff:
//------------------------

#2;
word <= 'hf3fffffffffffeff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1538
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6148: ir 'h%h !== 'hf", ir); end	// Vector No: 1537
assert (op === 'hff) else begin fail = 1; $display("Error 6149: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6150: extop 'h%h !== 0", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 6151: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// f3fffffffffffeff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffeff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1539
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6152: ir 'h%h !== 'hb", ir); end	// Vector No: 1538
assert (op === 'hf8) else begin fail = 1; $display("Error 6153: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6154: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6155: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffeff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffeff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1540
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6156: ir 'h%h !== 'hf", ir); end	// Vector No: 1539
assert (op === 'hf8) else begin fail = 1; $display("Error 6157: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6158: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6159: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffdff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffdff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1541
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6160: ir 'h%h !== 'hf", ir); end	// Vector No: 1540
assert (op === 'hff) else begin fail = 1; $display("Error 6161: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6162: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6163: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffdff:0:1:f:ff:1:ffdff:
//------------------------

#2;
word <= 'hfffffffff3fffdff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1542
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6164: ir 'h%h !== 'hf", ir); end	// Vector No: 1541
assert (op === 'hff) else begin fail = 1; $display("Error 6165: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6166: extop 'h%h !== 1", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 6167: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// fffffffff3fffdff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffdff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1543
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6168: ir 'h%h !== 'hf", ir); end	// Vector No: 1542
assert (op === 'hf8) else begin fail = 1; $display("Error 6169: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6170: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6171: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffdff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffdff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1544
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6172: ir 'h%h !== 'hf", ir); end	// Vector No: 1543
assert (op === 'hf0) else begin fail = 1; $display("Error 6173: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6174: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6175: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffdff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffdff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1545
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6176: ir 'h%h !== 'hf", ir); end	// Vector No: 1544
assert (op === 'hff) else begin fail = 1; $display("Error 6177: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6178: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6179: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffdff:0:1:f:ff:0:ffdff:
//------------------------

#2;
word <= 'hf3fffffffffffdff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1546
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6180: ir 'h%h !== 'hf", ir); end	// Vector No: 1545
assert (op === 'hff) else begin fail = 1; $display("Error 6181: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6182: extop 'h%h !== 0", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 6183: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// f3fffffffffffdff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffdff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1547
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6184: ir 'h%h !== 'hb", ir); end	// Vector No: 1546
assert (op === 'hf8) else begin fail = 1; $display("Error 6185: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6186: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6187: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffdff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffdff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1548
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6188: ir 'h%h !== 'hf", ir); end	// Vector No: 1547
assert (op === 'hf8) else begin fail = 1; $display("Error 6189: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6190: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6191: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffbff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fffbff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1549
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6192: ir 'h%h !== 'hf", ir); end	// Vector No: 1548
assert (op === 'hff) else begin fail = 1; $display("Error 6193: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6194: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6195: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fffbff:0:1:f:ff:1:ffbff:
//------------------------

#2;
word <= 'hfffffffff3fffbff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1550
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6196: ir 'h%h !== 'hf", ir); end	// Vector No: 1549
assert (op === 'hff) else begin fail = 1; $display("Error 6197: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6198: extop 'h%h !== 1", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 6199: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// fffffffff3fffbff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fffbff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1551
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6200: ir 'h%h !== 'hf", ir); end	// Vector No: 1550
assert (op === 'hf8) else begin fail = 1; $display("Error 6201: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6202: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6203: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fffbff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fffbff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1552
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6204: ir 'h%h !== 'hf", ir); end	// Vector No: 1551
assert (op === 'hf0) else begin fail = 1; $display("Error 6205: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6206: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6207: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffffbff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffffbff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1553
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6208: ir 'h%h !== 'hf", ir); end	// Vector No: 1552
assert (op === 'hff) else begin fail = 1; $display("Error 6209: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6210: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6211: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffffbff:0:1:f:ff:0:ffbff:
//------------------------

#2;
word <= 'hf3fffffffffffbff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1554
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6212: ir 'h%h !== 'hf", ir); end	// Vector No: 1553
assert (op === 'hff) else begin fail = 1; $display("Error 6213: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6214: extop 'h%h !== 0", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 6215: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// f3fffffffffffbff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffbff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1555
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6216: ir 'h%h !== 'hb", ir); end	// Vector No: 1554
assert (op === 'hf8) else begin fail = 1; $display("Error 6217: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6218: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6219: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffffbff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffffbff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1556
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6220: ir 'h%h !== 'hf", ir); end	// Vector No: 1555
assert (op === 'hf8) else begin fail = 1; $display("Error 6221: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6222: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6223: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fff7ff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fff7ff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1557
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6224: ir 'h%h !== 'hf", ir); end	// Vector No: 1556
assert (op === 'hff) else begin fail = 1; $display("Error 6225: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6226: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6227: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fff7ff:0:1:f:ff:1:ff7ff:
//------------------------

#2;
word <= 'hfffffffff3fff7ff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1558
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6228: ir 'h%h !== 'hf", ir); end	// Vector No: 1557
assert (op === 'hff) else begin fail = 1; $display("Error 6229: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6230: extop 'h%h !== 1", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 6231: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// fffffffff3fff7ff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fff7ff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1559
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6232: ir 'h%h !== 'hf", ir); end	// Vector No: 1558
assert (op === 'hf8) else begin fail = 1; $display("Error 6233: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6234: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6235: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fff7ff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3fff7ff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1560
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6236: ir 'h%h !== 'hf", ir); end	// Vector No: 1559
assert (op === 'hf0) else begin fail = 1; $display("Error 6237: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6238: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6239: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffffffff7ff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffff7ff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1561
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6240: ir 'h%h !== 'hf", ir); end	// Vector No: 1560
assert (op === 'hff) else begin fail = 1; $display("Error 6241: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6242: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6243: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffff7ff:0:1:f:ff:0:ff7ff:
//------------------------

#2;
word <= 'hf3fffffffffff7ff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1562
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6244: ir 'h%h !== 'hf", ir); end	// Vector No: 1561
assert (op === 'hff) else begin fail = 1; $display("Error 6245: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6246: extop 'h%h !== 0", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 6247: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// f3fffffffffff7ff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffff7ff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1563
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6248: ir 'h%h !== 'hb", ir); end	// Vector No: 1562
assert (op === 'hf8) else begin fail = 1; $display("Error 6249: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6250: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6251: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffff7ff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffff7ff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1564
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6252: ir 'h%h !== 'hf", ir); end	// Vector No: 1563
assert (op === 'hf8) else begin fail = 1; $display("Error 6253: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6254: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6255: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffefff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffefff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1565
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6256: ir 'h%h !== 'hf", ir); end	// Vector No: 1564
assert (op === 'hff) else begin fail = 1; $display("Error 6257: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6258: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6259: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffefff:0:1:f:fe:1:fefff:
//------------------------

#2;
word <= 'hfffffffff3ffefff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1566
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6260: ir 'h%h !== 'hf", ir); end	// Vector No: 1565
assert (op === 'hfe) else begin fail = 1; $display("Error 6261: op 'h%h !== 'hfe", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6262: extop 'h%h !== 1", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 6263: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// fffffffff3ffefff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffefff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1567
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6264: ir 'h%h !== 'hf", ir); end	// Vector No: 1566
assert (op === 'hf8) else begin fail = 1; $display("Error 6265: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6266: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6267: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffefff:1:1:f:f0:0:03ffe:
//------------------------

#2;
word <= 'hfffffffff3ffefff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1568
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6268: ir 'h%h !== 'hf", ir); end	// Vector No: 1567
assert (op === 'hf0) else begin fail = 1; $display("Error 6269: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6270: extop 'h%h !== 0", extop); end
assert (addr === 'h03ffe) else begin fail = 1; $display("Error 6271: addr 'h%h !== 'h03ffe", addr); end
#2;
clk <= 0;

// f3ffffffffffefff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffefff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1569
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6272: ir 'h%h !== 'hf", ir); end	// Vector No: 1568
assert (op === 'hff) else begin fail = 1; $display("Error 6273: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6274: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6275: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffefff:0:1:f:ff:0:fefff:
//------------------------

#2;
word <= 'hf3ffffffffffefff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1570
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6276: ir 'h%h !== 'hf", ir); end	// Vector No: 1569
assert (op === 'hff) else begin fail = 1; $display("Error 6277: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6278: extop 'h%h !== 0", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 6279: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// f3ffffffffffefff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffefff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1571
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6280: ir 'h%h !== 'hb", ir); end	// Vector No: 1570
assert (op === 'hf8) else begin fail = 1; $display("Error 6281: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6282: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6283: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffefff:1:1:f:f8:0:07ffe:
//------------------------

#2;
word <= 'hf3ffffffffffefff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1572
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6284: ir 'h%h !== 'hf", ir); end	// Vector No: 1571
assert (op === 'hf8) else begin fail = 1; $display("Error 6285: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6286: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffe) else begin fail = 1; $display("Error 6287: addr 'h%h !== 'h07ffe", addr); end
#2;
clk <= 0;

// fffffffff3ffdfff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffdfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1573
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6288: ir 'h%h !== 'hf", ir); end	// Vector No: 1572
assert (op === 'hff) else begin fail = 1; $display("Error 6289: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6290: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6291: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffdfff:0:1:f:fd:1:fdfff:
//------------------------

#2;
word <= 'hfffffffff3ffdfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1574
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6292: ir 'h%h !== 'hf", ir); end	// Vector No: 1573
assert (op === 'hfd) else begin fail = 1; $display("Error 6293: op 'h%h !== 'hfd", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6294: extop 'h%h !== 1", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 6295: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// fffffffff3ffdfff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffdfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1575
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6296: ir 'h%h !== 'hf", ir); end	// Vector No: 1574
assert (op === 'hf8) else begin fail = 1; $display("Error 6297: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6298: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6299: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffdfff:1:1:f:f0:0:03ffd:
//------------------------

#2;
word <= 'hfffffffff3ffdfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1576
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6300: ir 'h%h !== 'hf", ir); end	// Vector No: 1575
assert (op === 'hf0) else begin fail = 1; $display("Error 6301: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6302: extop 'h%h !== 0", extop); end
assert (addr === 'h03ffd) else begin fail = 1; $display("Error 6303: addr 'h%h !== 'h03ffd", addr); end
#2;
clk <= 0;

// f3ffffffffffdfff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffdfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1577
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6304: ir 'h%h !== 'hf", ir); end	// Vector No: 1576
assert (op === 'hff) else begin fail = 1; $display("Error 6305: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6306: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6307: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffdfff:0:1:f:ff:0:fdfff:
//------------------------

#2;
word <= 'hf3ffffffffffdfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1578
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6308: ir 'h%h !== 'hf", ir); end	// Vector No: 1577
assert (op === 'hff) else begin fail = 1; $display("Error 6309: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6310: extop 'h%h !== 0", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 6311: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// f3ffffffffffdfff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffdfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1579
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6312: ir 'h%h !== 'hb", ir); end	// Vector No: 1578
assert (op === 'hf8) else begin fail = 1; $display("Error 6313: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6314: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6315: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffdfff:1:1:f:f8:0:07ffd:
//------------------------

#2;
word <= 'hf3ffffffffffdfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1580
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6316: ir 'h%h !== 'hf", ir); end	// Vector No: 1579
assert (op === 'hf8) else begin fail = 1; $display("Error 6317: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6318: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffd) else begin fail = 1; $display("Error 6319: addr 'h%h !== 'h07ffd", addr); end
#2;
clk <= 0;

// fffffffff3ffbfff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffbfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1581
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6320: ir 'h%h !== 'hf", ir); end	// Vector No: 1580
assert (op === 'hff) else begin fail = 1; $display("Error 6321: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6322: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6323: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffbfff:0:1:f:fb:1:fbfff:
//------------------------

#2;
word <= 'hfffffffff3ffbfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1582
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6324: ir 'h%h !== 'hf", ir); end	// Vector No: 1581
assert (op === 'hfb) else begin fail = 1; $display("Error 6325: op 'h%h !== 'hfb", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6326: extop 'h%h !== 1", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 6327: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// fffffffff3ffbfff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffbfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1583
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6328: ir 'h%h !== 'hf", ir); end	// Vector No: 1582
assert (op === 'hf8) else begin fail = 1; $display("Error 6329: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6330: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6331: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffbfff:1:1:f:f0:0:03ffb:
//------------------------

#2;
word <= 'hfffffffff3ffbfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1584
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6332: ir 'h%h !== 'hf", ir); end	// Vector No: 1583
assert (op === 'hf0) else begin fail = 1; $display("Error 6333: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6334: extop 'h%h !== 0", extop); end
assert (addr === 'h03ffb) else begin fail = 1; $display("Error 6335: addr 'h%h !== 'h03ffb", addr); end
#2;
clk <= 0;

// f3ffffffffffbfff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffbfff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1585
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6336: ir 'h%h !== 'hf", ir); end	// Vector No: 1584
assert (op === 'hff) else begin fail = 1; $display("Error 6337: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6338: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6339: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffbfff:0:1:f:ff:0:fbfff:
//------------------------

#2;
word <= 'hf3ffffffffffbfff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1586
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6340: ir 'h%h !== 'hf", ir); end	// Vector No: 1585
assert (op === 'hff) else begin fail = 1; $display("Error 6341: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6342: extop 'h%h !== 0", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 6343: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// f3ffffffffffbfff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffbfff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1587
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6344: ir 'h%h !== 'hb", ir); end	// Vector No: 1586
assert (op === 'hf8) else begin fail = 1; $display("Error 6345: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6346: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6347: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffbfff:1:1:f:f8:0:07ffb:
//------------------------

#2;
word <= 'hf3ffffffffffbfff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1588
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6348: ir 'h%h !== 'hf", ir); end	// Vector No: 1587
assert (op === 'hf8) else begin fail = 1; $display("Error 6349: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6350: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffb) else begin fail = 1; $display("Error 6351: addr 'h%h !== 'h07ffb", addr); end
#2;
clk <= 0;

// fffffffff3ff7fff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ff7fff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1589
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6352: ir 'h%h !== 'hf", ir); end	// Vector No: 1588
assert (op === 'hff) else begin fail = 1; $display("Error 6353: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6354: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6355: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ff7fff:0:1:f:f7:1:f7fff:
//------------------------

#2;
word <= 'hfffffffff3ff7fff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1590
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6356: ir 'h%h !== 'hf", ir); end	// Vector No: 1589
assert (op === 'hf7) else begin fail = 1; $display("Error 6357: op 'h%h !== 'hf7", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6358: extop 'h%h !== 1", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 6359: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// fffffffff3ff7fff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ff7fff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1591
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6360: ir 'h%h !== 'hf", ir); end	// Vector No: 1590
assert (op === 'hf8) else begin fail = 1; $display("Error 6361: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6362: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6363: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ff7fff:1:1:f:f0:0:03ff7:
//------------------------

#2;
word <= 'hfffffffff3ff7fff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1592
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6364: ir 'h%h !== 'hf", ir); end	// Vector No: 1591
assert (op === 'hf0) else begin fail = 1; $display("Error 6365: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6366: extop 'h%h !== 0", extop); end
assert (addr === 'h03ff7) else begin fail = 1; $display("Error 6367: addr 'h%h !== 'h03ff7", addr); end
#2;
clk <= 0;

// f3ffffffffff7fff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffff7fff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1593
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6368: ir 'h%h !== 'hf", ir); end	// Vector No: 1592
assert (op === 'hff) else begin fail = 1; $display("Error 6369: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6370: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6371: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffff7fff:0:1:f:ff:0:f7fff:
//------------------------

#2;
word <= 'hf3ffffffffff7fff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1594
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6372: ir 'h%h !== 'hf", ir); end	// Vector No: 1593
assert (op === 'hff) else begin fail = 1; $display("Error 6373: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6374: extop 'h%h !== 0", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 6375: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// f3ffffffffff7fff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffff7fff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1595
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6376: ir 'h%h !== 'hb", ir); end	// Vector No: 1594
assert (op === 'hf8) else begin fail = 1; $display("Error 6377: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6378: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6379: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffff7fff:1:1:f:f8:0:07ff7:
//------------------------

#2;
word <= 'hf3ffffffffff7fff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1596
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6380: ir 'h%h !== 'hf", ir); end	// Vector No: 1595
assert (op === 'hf8) else begin fail = 1; $display("Error 6381: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6382: extop 'h%h !== 0", extop); end
assert (addr === 'h07ff7) else begin fail = 1; $display("Error 6383: addr 'h%h !== 'h07ff7", addr); end
#2;
clk <= 0;

// fffffffff3feffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3feffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1597
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6384: ir 'h%h !== 'hf", ir); end	// Vector No: 1596
assert (op === 'hff) else begin fail = 1; $display("Error 6385: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6386: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6387: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3feffff:0:1:f:ef:1:effff:
//------------------------

#2;
word <= 'hfffffffff3feffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1598
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6388: ir 'h%h !== 'hf", ir); end	// Vector No: 1597
assert (op === 'hef) else begin fail = 1; $display("Error 6389: op 'h%h !== 'hef", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6390: extop 'h%h !== 1", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 6391: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// fffffffff3feffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3feffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1599
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6392: ir 'h%h !== 'hf", ir); end	// Vector No: 1598
assert (op === 'hf8) else begin fail = 1; $display("Error 6393: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6394: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6395: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3feffff:1:1:f:f0:0:03fef:
//------------------------

#2;
word <= 'hfffffffff3feffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1600
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6396: ir 'h%h !== 'hf", ir); end	// Vector No: 1599
assert (op === 'hf0) else begin fail = 1; $display("Error 6397: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6398: extop 'h%h !== 0", extop); end
assert (addr === 'h03fef) else begin fail = 1; $display("Error 6399: addr 'h%h !== 'h03fef", addr); end
#2;
clk <= 0;

// f3fffffffffeffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffeffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1601
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6400: ir 'h%h !== 'hf", ir); end	// Vector No: 1600
assert (op === 'hff) else begin fail = 1; $display("Error 6401: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6402: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6403: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffeffff:0:1:f:ff:0:effff:
//------------------------

#2;
word <= 'hf3fffffffffeffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1602
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6404: ir 'h%h !== 'hf", ir); end	// Vector No: 1601
assert (op === 'hff) else begin fail = 1; $display("Error 6405: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6406: extop 'h%h !== 0", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 6407: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// f3fffffffffeffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffeffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1603
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6408: ir 'h%h !== 'hb", ir); end	// Vector No: 1602
assert (op === 'hf8) else begin fail = 1; $display("Error 6409: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6410: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6411: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffeffff:1:1:f:f8:0:07fef:
//------------------------

#2;
word <= 'hf3fffffffffeffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1604
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6412: ir 'h%h !== 'hf", ir); end	// Vector No: 1603
assert (op === 'hf8) else begin fail = 1; $display("Error 6413: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6414: extop 'h%h !== 0", extop); end
assert (addr === 'h07fef) else begin fail = 1; $display("Error 6415: addr 'h%h !== 'h07fef", addr); end
#2;
clk <= 0;

// fffffffff3fdffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fdffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1605
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6416: ir 'h%h !== 'hf", ir); end	// Vector No: 1604
assert (op === 'hff) else begin fail = 1; $display("Error 6417: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6418: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6419: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fdffff:0:1:f:df:1:dffff:
//------------------------

#2;
word <= 'hfffffffff3fdffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1606
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6420: ir 'h%h !== 'hf", ir); end	// Vector No: 1605
assert (op === 'hdf) else begin fail = 1; $display("Error 6421: op 'h%h !== 'hdf", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6422: extop 'h%h !== 1", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 6423: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// fffffffff3fdffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fdffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1607
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6424: ir 'h%h !== 'hf", ir); end	// Vector No: 1606
assert (op === 'hf8) else begin fail = 1; $display("Error 6425: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6426: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6427: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fdffff:1:1:f:f0:0:03fdf:
//------------------------

#2;
word <= 'hfffffffff3fdffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1608
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6428: ir 'h%h !== 'hf", ir); end	// Vector No: 1607
assert (op === 'hf0) else begin fail = 1; $display("Error 6429: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6430: extop 'h%h !== 0", extop); end
assert (addr === 'h03fdf) else begin fail = 1; $display("Error 6431: addr 'h%h !== 'h03fdf", addr); end
#2;
clk <= 0;

// f3fffffffffdffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffdffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1609
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6432: ir 'h%h !== 'hf", ir); end	// Vector No: 1608
assert (op === 'hff) else begin fail = 1; $display("Error 6433: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6434: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6435: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffdffff:0:1:f:ff:0:dffff:
//------------------------

#2;
word <= 'hf3fffffffffdffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1610
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6436: ir 'h%h !== 'hf", ir); end	// Vector No: 1609
assert (op === 'hff) else begin fail = 1; $display("Error 6437: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6438: extop 'h%h !== 0", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 6439: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// f3fffffffffdffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffdffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1611
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6440: ir 'h%h !== 'hb", ir); end	// Vector No: 1610
assert (op === 'hf8) else begin fail = 1; $display("Error 6441: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6442: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6443: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffdffff:1:1:f:f8:0:07fdf:
//------------------------

#2;
word <= 'hf3fffffffffdffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1612
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6444: ir 'h%h !== 'hf", ir); end	// Vector No: 1611
assert (op === 'hf8) else begin fail = 1; $display("Error 6445: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6446: extop 'h%h !== 0", extop); end
assert (addr === 'h07fdf) else begin fail = 1; $display("Error 6447: addr 'h%h !== 'h07fdf", addr); end
#2;
clk <= 0;

// fffffffff3fbffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3fbffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1613
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6448: ir 'h%h !== 'hf", ir); end	// Vector No: 1612
assert (op === 'hff) else begin fail = 1; $display("Error 6449: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6450: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6451: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3fbffff:0:1:f:bf:1:bffff:
//------------------------

#2;
word <= 'hfffffffff3fbffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1614
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6452: ir 'h%h !== 'hf", ir); end	// Vector No: 1613
assert (op === 'hbf) else begin fail = 1; $display("Error 6453: op 'h%h !== 'hbf", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6454: extop 'h%h !== 1", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 6455: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// fffffffff3fbffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3fbffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1615
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6456: ir 'h%h !== 'hf", ir); end	// Vector No: 1614
assert (op === 'hf8) else begin fail = 1; $display("Error 6457: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6458: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6459: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3fbffff:1:1:f:f0:0:03fbf:
//------------------------

#2;
word <= 'hfffffffff3fbffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1616
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6460: ir 'h%h !== 'hf", ir); end	// Vector No: 1615
assert (op === 'hf0) else begin fail = 1; $display("Error 6461: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6462: extop 'h%h !== 0", extop); end
assert (addr === 'h03fbf) else begin fail = 1; $display("Error 6463: addr 'h%h !== 'h03fbf", addr); end
#2;
clk <= 0;

// f3fffffffffbffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffffbffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1617
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6464: ir 'h%h !== 'hf", ir); end	// Vector No: 1616
assert (op === 'hff) else begin fail = 1; $display("Error 6465: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6466: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6467: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffffbffff:0:1:f:ff:0:bffff:
//------------------------

#2;
word <= 'hf3fffffffffbffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1618
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6468: ir 'h%h !== 'hf", ir); end	// Vector No: 1617
assert (op === 'hff) else begin fail = 1; $display("Error 6469: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6470: extop 'h%h !== 0", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 6471: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// f3fffffffffbffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffffbffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1619
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6472: ir 'h%h !== 'hb", ir); end	// Vector No: 1618
assert (op === 'hf8) else begin fail = 1; $display("Error 6473: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6474: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6475: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffffbffff:1:1:f:f8:0:07fbf:
//------------------------

#2;
word <= 'hf3fffffffffbffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1620
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6476: ir 'h%h !== 'hf", ir); end	// Vector No: 1619
assert (op === 'hf8) else begin fail = 1; $display("Error 6477: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6478: extop 'h%h !== 0", extop); end
assert (addr === 'h07fbf) else begin fail = 1; $display("Error 6479: addr 'h%h !== 'h07fbf", addr); end
#2;
clk <= 0;

// fffffffff3f7ffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3f7ffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1621
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6480: ir 'h%h !== 'hf", ir); end	// Vector No: 1620
assert (op === 'hff) else begin fail = 1; $display("Error 6481: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6482: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6483: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3f7ffff:0:1:f:7f:1:7ffff:
//------------------------

#2;
word <= 'hfffffffff3f7ffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1622
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6484: ir 'h%h !== 'hf", ir); end	// Vector No: 1621
assert (op === 'h7f) else begin fail = 1; $display("Error 6485: op 'h%h !== 'h7f", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6486: extop 'h%h !== 1", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 6487: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// fffffffff3f7ffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3f7ffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1623
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6488: ir 'h%h !== 'hf", ir); end	// Vector No: 1622
assert (op === 'hf8) else begin fail = 1; $display("Error 6489: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6490: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6491: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3f7ffff:1:1:f:f0:0:03f7f:
//------------------------

#2;
word <= 'hfffffffff3f7ffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1624
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6492: ir 'h%h !== 'hf", ir); end	// Vector No: 1623
assert (op === 'hf0) else begin fail = 1; $display("Error 6493: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6494: extop 'h%h !== 0", extop); end
assert (addr === 'h03f7f) else begin fail = 1; $display("Error 6495: addr 'h%h !== 'h03f7f", addr); end
#2;
clk <= 0;

// f3fffffffff7ffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffff7ffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1625
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6496: ir 'h%h !== 'hf", ir); end	// Vector No: 1624
assert (op === 'hff) else begin fail = 1; $display("Error 6497: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6498: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6499: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffff7ffff:0:1:f:ff:0:7ffff:
//------------------------

#2;
word <= 'hf3fffffffff7ffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1626
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6500: ir 'h%h !== 'hf", ir); end	// Vector No: 1625
assert (op === 'hff) else begin fail = 1; $display("Error 6501: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6502: extop 'h%h !== 0", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 6503: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// f3fffffffff7ffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffff7ffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1627
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6504: ir 'h%h !== 'hb", ir); end	// Vector No: 1626
assert (op === 'hf8) else begin fail = 1; $display("Error 6505: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6506: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6507: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffff7ffff:1:1:f:f8:0:07f7f:
//------------------------

#2;
word <= 'hf3fffffffff7ffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1628
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6508: ir 'h%h !== 'hf", ir); end	// Vector No: 1627
assert (op === 'hf8) else begin fail = 1; $display("Error 6509: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6510: extop 'h%h !== 0", extop); end
assert (addr === 'h07f7f) else begin fail = 1; $display("Error 6511: addr 'h%h !== 'h07f7f", addr); end
#2;
clk <= 0;

// fffffffff3ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1629
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6512: ir 'h%h !== 'hf", ir); end	// Vector No: 1628
assert (op === 'hff) else begin fail = 1; $display("Error 6513: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6514: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6515: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1630
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6516: ir 'h%h !== 'hf", ir); end	// Vector No: 1629
assert (op === 'hff) else begin fail = 1; $display("Error 6517: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6518: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6519: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffff3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1631
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6520: ir 'h%h !== 'hf", ir); end	// Vector No: 1630
assert (op === 'hf8) else begin fail = 1; $display("Error 6521: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6522: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6523: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1632
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6524: ir 'h%h !== 'hf", ir); end	// Vector No: 1631
assert (op === 'hf0) else begin fail = 1; $display("Error 6525: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6526: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6527: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffefffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffefffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1633
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6528: ir 'h%h !== 'hf", ir); end	// Vector No: 1632
assert (op === 'hff) else begin fail = 1; $display("Error 6529: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6530: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6531: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffefffff:0:1:f:fe:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffffefffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1634
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6532: ir 'h%h !== 'hf", ir); end	// Vector No: 1633
assert (op === 'hfe) else begin fail = 1; $display("Error 6533: op 'h%h !== 'hfe", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6534: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6535: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffefffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffefffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1635
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6536: ir 'h%h !== 'hb", ir); end	// Vector No: 1634
assert (op === 'hf8) else begin fail = 1; $display("Error 6537: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6538: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6539: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffefffff:1:1:f:f8:0:07eff:
//------------------------

#2;
word <= 'hf3ffffffffefffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1636
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6540: ir 'h%h !== 'hf", ir); end	// Vector No: 1635
assert (op === 'hf8) else begin fail = 1; $display("Error 6541: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6542: extop 'h%h !== 0", extop); end
assert (addr === 'h07eff) else begin fail = 1; $display("Error 6543: addr 'h%h !== 'h07eff", addr); end
#2;
clk <= 0;

// f3ffffffffdfffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffdfffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1637
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6544: ir 'h%h !== 'hf", ir); end	// Vector No: 1636
assert (op === 'hff) else begin fail = 1; $display("Error 6545: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6546: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6547: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffdfffff:0:1:f:fd:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffffdfffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1638
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6548: ir 'h%h !== 'hf", ir); end	// Vector No: 1637
assert (op === 'hfd) else begin fail = 1; $display("Error 6549: op 'h%h !== 'hfd", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6550: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6551: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffdfffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffdfffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1639
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6552: ir 'h%h !== 'hb", ir); end	// Vector No: 1638
assert (op === 'hf8) else begin fail = 1; $display("Error 6553: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6554: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6555: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffdfffff:1:1:f:f8:0:07dff:
//------------------------

#2;
word <= 'hf3ffffffffdfffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1640
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6556: ir 'h%h !== 'hf", ir); end	// Vector No: 1639
assert (op === 'hf8) else begin fail = 1; $display("Error 6557: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6558: extop 'h%h !== 0", extop); end
assert (addr === 'h07dff) else begin fail = 1; $display("Error 6559: addr 'h%h !== 'h07dff", addr); end
#2;
clk <= 0;

// f3ffffffffbfffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffbfffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1641
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6560: ir 'h%h !== 'hf", ir); end	// Vector No: 1640
assert (op === 'hff) else begin fail = 1; $display("Error 6561: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6562: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6563: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffbfffff:0:1:f:fb:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffffbfffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1642
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6564: ir 'h%h !== 'hf", ir); end	// Vector No: 1641
assert (op === 'hfb) else begin fail = 1; $display("Error 6565: op 'h%h !== 'hfb", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6566: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6567: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffbfffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffbfffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1643
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6568: ir 'h%h !== 'hb", ir); end	// Vector No: 1642
assert (op === 'hf8) else begin fail = 1; $display("Error 6569: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6570: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6571: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffbfffff:1:1:f:f8:0:07bff:
//------------------------

#2;
word <= 'hf3ffffffffbfffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1644
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6572: ir 'h%h !== 'hf", ir); end	// Vector No: 1643
assert (op === 'hf8) else begin fail = 1; $display("Error 6573: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6574: extop 'h%h !== 0", extop); end
assert (addr === 'h07bff) else begin fail = 1; $display("Error 6575: addr 'h%h !== 'h07bff", addr); end
#2;
clk <= 0;

// f3ffffffff7fffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffff7fffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1645
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6576: ir 'h%h !== 'hf", ir); end	// Vector No: 1644
assert (op === 'hff) else begin fail = 1; $display("Error 6577: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6578: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6579: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffff7fffff:0:1:f:f7:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffff7fffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1646
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6580: ir 'h%h !== 'hf", ir); end	// Vector No: 1645
assert (op === 'hf7) else begin fail = 1; $display("Error 6581: op 'h%h !== 'hf7", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6582: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6583: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffff7fffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffff7fffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1647
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6584: ir 'h%h !== 'hb", ir); end	// Vector No: 1646
assert (op === 'hf8) else begin fail = 1; $display("Error 6585: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6586: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6587: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffff7fffff:1:1:f:f8:0:077ff:
//------------------------

#2;
word <= 'hf3ffffffff7fffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1648
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6588: ir 'h%h !== 'hf", ir); end	// Vector No: 1647
assert (op === 'hf8) else begin fail = 1; $display("Error 6589: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6590: extop 'h%h !== 0", extop); end
assert (addr === 'h077ff) else begin fail = 1; $display("Error 6591: addr 'h%h !== 'h077ff", addr); end
#2;
clk <= 0;

// f3fffffffeffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffeffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1649
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6592: ir 'h%h !== 'hf", ir); end	// Vector No: 1648
assert (op === 'hff) else begin fail = 1; $display("Error 6593: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6594: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6595: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffeffffff:0:1:f:ef:0:fffff:
//------------------------

#2;
word <= 'hf3fffffffeffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1650
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6596: ir 'h%h !== 'hf", ir); end	// Vector No: 1649
assert (op === 'hef) else begin fail = 1; $display("Error 6597: op 'h%h !== 'hef", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6598: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6599: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffeffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffeffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1651
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6600: ir 'h%h !== 'hb", ir); end	// Vector No: 1650
assert (op === 'hf8) else begin fail = 1; $display("Error 6601: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6602: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6603: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffeffffff:1:1:f:f8:0:06fff:
//------------------------

#2;
word <= 'hf3fffffffeffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1652
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6604: ir 'h%h !== 'hf", ir); end	// Vector No: 1651
assert (op === 'hf8) else begin fail = 1; $display("Error 6605: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6606: extop 'h%h !== 0", extop); end
assert (addr === 'h06fff) else begin fail = 1; $display("Error 6607: addr 'h%h !== 'h06fff", addr); end
#2;
clk <= 0;

// f3fffffffdffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffdffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1653
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6608: ir 'h%h !== 'hf", ir); end	// Vector No: 1652
assert (op === 'hff) else begin fail = 1; $display("Error 6609: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6610: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6611: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffdffffff:0:1:f:df:0:fffff:
//------------------------

#2;
word <= 'hf3fffffffdffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1654
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6612: ir 'h%h !== 'hf", ir); end	// Vector No: 1653
assert (op === 'hdf) else begin fail = 1; $display("Error 6613: op 'h%h !== 'hdf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6614: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6615: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffdffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffdffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1655
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6616: ir 'h%h !== 'hb", ir); end	// Vector No: 1654
assert (op === 'hf8) else begin fail = 1; $display("Error 6617: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6618: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6619: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffdffffff:1:1:f:f8:0:05fff:
//------------------------

#2;
word <= 'hf3fffffffdffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1656
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6620: ir 'h%h !== 'hf", ir); end	// Vector No: 1655
assert (op === 'hf8) else begin fail = 1; $display("Error 6621: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6622: extop 'h%h !== 0", extop); end
assert (addr === 'h05fff) else begin fail = 1; $display("Error 6623: addr 'h%h !== 'h05fff", addr); end
#2;
clk <= 0;

// f3fffffffbffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffffbffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1657
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6624: ir 'h%h !== 'hf", ir); end	// Vector No: 1656
assert (op === 'hff) else begin fail = 1; $display("Error 6625: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6626: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6627: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffbffffff:0:1:f:bf:0:fffff:
//------------------------

#2;
word <= 'hf3fffffffbffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1658
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6628: ir 'h%h !== 'hf", ir); end	// Vector No: 1657
assert (op === 'hbf) else begin fail = 1; $display("Error 6629: op 'h%h !== 'hbf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6630: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6631: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffffbffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffffbffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1659
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6632: ir 'h%h !== 'hb", ir); end	// Vector No: 1658
assert (op === 'hf8) else begin fail = 1; $display("Error 6633: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6634: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6635: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffffbffffff:1:1:f:f8:0:03fff:
//------------------------

#2;
word <= 'hf3fffffffbffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1660
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6636: ir 'h%h !== 'hf", ir); end	// Vector No: 1659
assert (op === 'hf8) else begin fail = 1; $display("Error 6637: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6638: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6639: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffff7ffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3fffffff7ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1661
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6640: ir 'h%h !== 'hf", ir); end	// Vector No: 1660
assert (op === 'hff) else begin fail = 1; $display("Error 6641: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6642: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6643: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffff7ffffff:0:1:f:7f:0:fffff:
//------------------------

#2;
word <= 'hf3fffffff7ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1662
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6644: ir 'h%h !== 'hf", ir); end	// Vector No: 1661
assert (op === 'h7f) else begin fail = 1; $display("Error 6645: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6646: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6647: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffff7ffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffff7ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1663
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6648: ir 'h%h !== 'hb", ir); end	// Vector No: 1662
assert (op === 'hf8) else begin fail = 1; $display("Error 6649: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6650: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6651: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffff7ffffff:1:1:f:f0:0:07fff:
//------------------------

#2;
word <= 'hf3fffffff7ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1664
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6652: ir 'h%h !== 'hf", ir); end	// Vector No: 1663
assert (op === 'hf0) else begin fail = 1; $display("Error 6653: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6654: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6655: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffe3ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffe3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1665
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6656: ir 'h%h !== 'hf", ir); end	// Vector No: 1664
assert (op === 'hff) else begin fail = 1; $display("Error 6657: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6658: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6659: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffe3ffffff:0:1:e:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffffe3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1666
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 6660: ir 'h%h !== 'he", ir); end	// Vector No: 1665
assert (op === 'hff) else begin fail = 1; $display("Error 6661: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6662: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6663: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffe3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffe3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1667
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6664: ir 'h%h !== 'hf", ir); end	// Vector No: 1666
assert (op === 'hf8) else begin fail = 1; $display("Error 6665: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6666: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6667: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffe3ffffff:1:1:f:e0:0:03fff:
//------------------------

#2;
word <= 'hffffffffe3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1668
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6668: ir 'h%h !== 'hf", ir); end	// Vector No: 1667
assert (op === 'he0) else begin fail = 1; $display("Error 6669: op 'h%h !== 'he0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6670: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6671: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffefffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffefffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1669
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6672: ir 'h%h !== 'hf", ir); end	// Vector No: 1668
assert (op === 'hff) else begin fail = 1; $display("Error 6673: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6674: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6675: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffefffffff:0:1:e:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffefffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1670
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 6676: ir 'h%h !== 'he", ir); end	// Vector No: 1669
assert (op === 'hff) else begin fail = 1; $display("Error 6677: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6678: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6679: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffefffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffefffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1671
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6680: ir 'h%h !== 'hb", ir); end	// Vector No: 1670
assert (op === 'hf8) else begin fail = 1; $display("Error 6681: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6682: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6683: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffefffffff:1:1:f:e8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffefffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1672
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6684: ir 'h%h !== 'hf", ir); end	// Vector No: 1671
assert (op === 'he8) else begin fail = 1; $display("Error 6685: op 'h%h !== 'he8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6686: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6687: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffd3ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffd3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1673
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6688: ir 'h%h !== 'hf", ir); end	// Vector No: 1672
assert (op === 'hff) else begin fail = 1; $display("Error 6689: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6690: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6691: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffd3ffffff:0:1:d:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffffd3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1674
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 6692: ir 'h%h !== 'hd", ir); end	// Vector No: 1673
assert (op === 'hff) else begin fail = 1; $display("Error 6693: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6694: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6695: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffd3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffd3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1675
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6696: ir 'h%h !== 'hf", ir); end	// Vector No: 1674
assert (op === 'hf8) else begin fail = 1; $display("Error 6697: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6698: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6699: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffd3ffffff:1:1:f:d0:0:03fff:
//------------------------

#2;
word <= 'hffffffffd3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1676
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6700: ir 'h%h !== 'hf", ir); end	// Vector No: 1675
assert (op === 'hd0) else begin fail = 1; $display("Error 6701: op 'h%h !== 'hd0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6702: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6703: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffdfffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffdfffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1677
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6704: ir 'h%h !== 'hf", ir); end	// Vector No: 1676
assert (op === 'hff) else begin fail = 1; $display("Error 6705: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6706: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6707: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffdfffffff:0:1:d:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffdfffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1678
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 6708: ir 'h%h !== 'hd", ir); end	// Vector No: 1677
assert (op === 'hff) else begin fail = 1; $display("Error 6709: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6710: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6711: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffdfffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffdfffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1679
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6712: ir 'h%h !== 'hb", ir); end	// Vector No: 1678
assert (op === 'hf8) else begin fail = 1; $display("Error 6713: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6714: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6715: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffdfffffff:1:1:f:d8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffdfffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1680
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6716: ir 'h%h !== 'hf", ir); end	// Vector No: 1679
assert (op === 'hd8) else begin fail = 1; $display("Error 6717: op 'h%h !== 'hd8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6718: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6719: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffb3ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffffb3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1681
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6720: ir 'h%h !== 'hf", ir); end	// Vector No: 1680
assert (op === 'hff) else begin fail = 1; $display("Error 6721: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6722: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6723: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffb3ffffff:0:1:b:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffffb3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1682
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6724: ir 'h%h !== 'hb", ir); end	// Vector No: 1681
assert (op === 'hff) else begin fail = 1; $display("Error 6725: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6726: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6727: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffffb3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffffb3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1683
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6728: ir 'h%h !== 'hf", ir); end	// Vector No: 1682
assert (op === 'hf8) else begin fail = 1; $display("Error 6729: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6730: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6731: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffffb3ffffff:1:1:f:b0:0:03fff:
//------------------------

#2;
word <= 'hffffffffb3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1684
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6732: ir 'h%h !== 'hf", ir); end	// Vector No: 1683
assert (op === 'hb0) else begin fail = 1; $display("Error 6733: op 'h%h !== 'hb0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6734: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6735: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffbfffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffbfffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1685
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6736: ir 'h%h !== 'hf", ir); end	// Vector No: 1684
assert (op === 'hff) else begin fail = 1; $display("Error 6737: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6738: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6739: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffbfffffff:0:1:b:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffbfffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1686
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6740: ir 'h%h !== 'hb", ir); end	// Vector No: 1685
assert (op === 'hff) else begin fail = 1; $display("Error 6741: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6742: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6743: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffbfffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffbfffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1687
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6744: ir 'h%h !== 'hb", ir); end	// Vector No: 1686
assert (op === 'hf8) else begin fail = 1; $display("Error 6745: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6746: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6747: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffbfffffff:1:1:f:b8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffbfffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1688
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6748: ir 'h%h !== 'hf", ir); end	// Vector No: 1687
assert (op === 'hb8) else begin fail = 1; $display("Error 6749: op 'h%h !== 'hb8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6750: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6751: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffff73ffffff:0:0:f:ff:0:fffff:
//------------------------

#2;
word <= 'hffffffff73ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1689
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6752: ir 'h%h !== 'hf", ir); end	// Vector No: 1688
assert (op === 'hff) else begin fail = 1; $display("Error 6753: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6754: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6755: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffff73ffffff:0:1:7:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffff73ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1690
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 6756: ir 'h%h !== 'h7", ir); end	// Vector No: 1689
assert (op === 'hff) else begin fail = 1; $display("Error 6757: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6758: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6759: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffff73ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hffffffff73ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1691
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6760: ir 'h%h !== 'hf", ir); end	// Vector No: 1690
assert (op === 'hf8) else begin fail = 1; $display("Error 6761: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6762: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6763: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffff73ffffff:1:1:f:73:0:07fff:
//------------------------

#2;
word <= 'hffffffff73ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1692
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6764: ir 'h%h !== 'hf", ir); end	// Vector No: 1691
assert (op === 'h73) else begin fail = 1; $display("Error 6765: op 'h%h !== 'h73", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6766: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6767: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffff7fffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffff7fffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1693
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6768: ir 'h%h !== 'hf", ir); end	// Vector No: 1692
assert (op === 'hff) else begin fail = 1; $display("Error 6769: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6770: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6771: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffff7fffffff:0:1:7:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffff7fffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1694
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 6772: ir 'h%h !== 'h7", ir); end	// Vector No: 1693
assert (op === 'hff) else begin fail = 1; $display("Error 6773: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6774: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6775: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffff7fffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffff7fffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1695
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6776: ir 'h%h !== 'hb", ir); end	// Vector No: 1694
assert (op === 'hf8) else begin fail = 1; $display("Error 6777: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6778: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6779: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffff7fffffff:1:1:f:7f:0:07fff:
//------------------------

#2;
word <= 'hf3ffffff7fffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1696
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6780: ir 'h%h !== 'hf", ir); end	// Vector No: 1695
assert (op === 'h7f) else begin fail = 1; $display("Error 6781: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6782: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6783: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffef3ffffff:0:0:f:ff:0:ffffe:
//------------------------

#2;
word <= 'hfffffffef3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1697
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6784: ir 'h%h !== 'hf", ir); end	// Vector No: 1696
assert (op === 'hff) else begin fail = 1; $display("Error 6785: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6786: extop 'h%h !== 0", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 6787: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// fffffffef3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffffef3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1698
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6788: ir 'h%h !== 'hf", ir); end	// Vector No: 1697
assert (op === 'hff) else begin fail = 1; $display("Error 6789: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6790: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6791: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffef3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffef3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1699
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6792: ir 'h%h !== 'hf", ir); end	// Vector No: 1698
assert (op === 'hf8) else begin fail = 1; $display("Error 6793: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6794: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6795: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffef3ffffff:1:1:e:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffef3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1700
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 6796: ir 'h%h !== 'he", ir); end	// Vector No: 1699
assert (op === 'hf0) else begin fail = 1; $display("Error 6797: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6798: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6799: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffeffffffff:0:0:f:ff:1:ffffe:
//------------------------

#2;
word <= 'hf3fffffeffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1701
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6800: ir 'h%h !== 'hf", ir); end	// Vector No: 1700
assert (op === 'hff) else begin fail = 1; $display("Error 6801: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6802: extop 'h%h !== 1", extop); end
assert (addr === 'hffffe) else begin fail = 1; $display("Error 6803: addr 'h%h !== 'hffffe", addr); end
#2;
clk <= 0;

// f3fffffeffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffffeffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1702
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6804: ir 'h%h !== 'hf", ir); end	// Vector No: 1701
assert (op === 'hff) else begin fail = 1; $display("Error 6805: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6806: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6807: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffeffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffeffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1703
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6808: ir 'h%h !== 'hb", ir); end	// Vector No: 1702
assert (op === 'hf8) else begin fail = 1; $display("Error 6809: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6810: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6811: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffeffffffff:1:1:e:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffeffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1704
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 6812: ir 'h%h !== 'he", ir); end	// Vector No: 1703
assert (op === 'hf8) else begin fail = 1; $display("Error 6813: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6814: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6815: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffdf3ffffff:0:0:f:ff:0:ffffd:
//------------------------

#2;
word <= 'hfffffffdf3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1705
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6816: ir 'h%h !== 'hf", ir); end	// Vector No: 1704
assert (op === 'hff) else begin fail = 1; $display("Error 6817: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6818: extop 'h%h !== 0", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 6819: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// fffffffdf3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffffdf3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1706
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6820: ir 'h%h !== 'hf", ir); end	// Vector No: 1705
assert (op === 'hff) else begin fail = 1; $display("Error 6821: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6822: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6823: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffdf3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffdf3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1707
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6824: ir 'h%h !== 'hf", ir); end	// Vector No: 1706
assert (op === 'hf8) else begin fail = 1; $display("Error 6825: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6826: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6827: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffdf3ffffff:1:1:d:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffdf3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1708
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 6828: ir 'h%h !== 'hd", ir); end	// Vector No: 1707
assert (op === 'hf0) else begin fail = 1; $display("Error 6829: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6830: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6831: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffdffffffff:0:0:f:ff:1:ffffd:
//------------------------

#2;
word <= 'hf3fffffdffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1709
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6832: ir 'h%h !== 'hf", ir); end	// Vector No: 1708
assert (op === 'hff) else begin fail = 1; $display("Error 6833: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6834: extop 'h%h !== 1", extop); end
assert (addr === 'hffffd) else begin fail = 1; $display("Error 6835: addr 'h%h !== 'hffffd", addr); end
#2;
clk <= 0;

// f3fffffdffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffffdffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1710
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6836: ir 'h%h !== 'hf", ir); end	// Vector No: 1709
assert (op === 'hff) else begin fail = 1; $display("Error 6837: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6838: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6839: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffdffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffdffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1711
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6840: ir 'h%h !== 'hb", ir); end	// Vector No: 1710
assert (op === 'hf8) else begin fail = 1; $display("Error 6841: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6842: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6843: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffdffffffff:1:1:d:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffdffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1712
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 6844: ir 'h%h !== 'hd", ir); end	// Vector No: 1711
assert (op === 'hf8) else begin fail = 1; $display("Error 6845: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6846: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6847: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffbf3ffffff:0:0:f:ff:0:ffffb:
//------------------------

#2;
word <= 'hfffffffbf3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1713
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6848: ir 'h%h !== 'hf", ir); end	// Vector No: 1712
assert (op === 'hff) else begin fail = 1; $display("Error 6849: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6850: extop 'h%h !== 0", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 6851: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// fffffffbf3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffffbf3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1714
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6852: ir 'h%h !== 'hf", ir); end	// Vector No: 1713
assert (op === 'hff) else begin fail = 1; $display("Error 6853: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6854: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6855: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffffbf3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffffbf3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1715
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6856: ir 'h%h !== 'hf", ir); end	// Vector No: 1714
assert (op === 'hf8) else begin fail = 1; $display("Error 6857: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6858: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6859: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffffbf3ffffff:1:1:b:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffffbf3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1716
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6860: ir 'h%h !== 'hb", ir); end	// Vector No: 1715
assert (op === 'hf0) else begin fail = 1; $display("Error 6861: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6862: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6863: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffffbffffffff:0:0:f:ff:1:ffffb:
//------------------------

#2;
word <= 'hf3fffffbffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1717
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6864: ir 'h%h !== 'hf", ir); end	// Vector No: 1716
assert (op === 'hff) else begin fail = 1; $display("Error 6865: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6866: extop 'h%h !== 1", extop); end
assert (addr === 'hffffb) else begin fail = 1; $display("Error 6867: addr 'h%h !== 'hffffb", addr); end
#2;
clk <= 0;

// f3fffffbffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffffbffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1718
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6868: ir 'h%h !== 'hf", ir); end	// Vector No: 1717
assert (op === 'hff) else begin fail = 1; $display("Error 6869: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6870: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6871: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffffbffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffbffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1719
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6872: ir 'h%h !== 'hb", ir); end	// Vector No: 1718
assert (op === 'hf8) else begin fail = 1; $display("Error 6873: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6874: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6875: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffffbffffffff:1:1:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffffbffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1720
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6876: ir 'h%h !== 'hb", ir); end	// Vector No: 1719
assert (op === 'hf8) else begin fail = 1; $display("Error 6877: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6878: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6879: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffff7f3ffffff:0:0:f:ff:0:ffff7:
//------------------------

#2;
word <= 'hfffffff7f3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1721
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6880: ir 'h%h !== 'hf", ir); end	// Vector No: 1720
assert (op === 'hff) else begin fail = 1; $display("Error 6881: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6882: extop 'h%h !== 0", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 6883: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// fffffff7f3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffff7f3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1722
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6884: ir 'h%h !== 'hf", ir); end	// Vector No: 1721
assert (op === 'hff) else begin fail = 1; $display("Error 6885: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6886: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6887: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffff7f3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hfffffff7f3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1723
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6888: ir 'h%h !== 'hf", ir); end	// Vector No: 1722
assert (op === 'hf8) else begin fail = 1; $display("Error 6889: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6890: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6891: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffff7f3ffffff:1:1:7:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffff7f3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1724
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 6892: ir 'h%h !== 'h7", ir); end	// Vector No: 1723
assert (op === 'hf0) else begin fail = 1; $display("Error 6893: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6894: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6895: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffff7ffffffff:0:0:f:ff:1:ffff7:
//------------------------

#2;
word <= 'hf3fffff7ffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1725
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6896: ir 'h%h !== 'hf", ir); end	// Vector No: 1724
assert (op === 'hff) else begin fail = 1; $display("Error 6897: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6898: extop 'h%h !== 1", extop); end
assert (addr === 'hffff7) else begin fail = 1; $display("Error 6899: addr 'h%h !== 'hffff7", addr); end
#2;
clk <= 0;

// f3fffff7ffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffff7ffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1726
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6900: ir 'h%h !== 'hf", ir); end	// Vector No: 1725
assert (op === 'hff) else begin fail = 1; $display("Error 6901: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6902: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6903: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffff7ffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffff7ffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1727
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6904: ir 'h%h !== 'hb", ir); end	// Vector No: 1726
assert (op === 'hf8) else begin fail = 1; $display("Error 6905: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6906: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6907: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3fffff7ffffffff:1:1:7:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffff7ffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1728
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 6908: ir 'h%h !== 'h7", ir); end	// Vector No: 1727
assert (op === 'hf8) else begin fail = 1; $display("Error 6909: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6910: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6911: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffeff3ffffff:0:0:f:ff:0:fffef:
//------------------------

#2;
word <= 'hffffffeff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1729
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6912: ir 'h%h !== 'hf", ir); end	// Vector No: 1728
assert (op === 'hff) else begin fail = 1; $display("Error 6913: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6914: extop 'h%h !== 0", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 6915: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// ffffffeff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffeff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1730
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6916: ir 'h%h !== 'hf", ir); end	// Vector No: 1729
assert (op === 'hff) else begin fail = 1; $display("Error 6917: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6918: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6919: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffeff3ffffff:1:0:f:f8:0:07ffe:
//------------------------

#2;
word <= 'hffffffeff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1731
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6920: ir 'h%h !== 'hf", ir); end	// Vector No: 1730
assert (op === 'hf8) else begin fail = 1; $display("Error 6921: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6922: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffe) else begin fail = 1; $display("Error 6923: addr 'h%h !== 'h07ffe", addr); end
#2;
clk <= 0;

// ffffffeff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffffeff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1732
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6924: ir 'h%h !== 'hf", ir); end	// Vector No: 1731
assert (op === 'hf0) else begin fail = 1; $display("Error 6925: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6926: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6927: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffefffffffff:0:0:f:ff:1:fffef:
//------------------------

#2;
word <= 'hf3ffffefffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1733
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6928: ir 'h%h !== 'hf", ir); end	// Vector No: 1732
assert (op === 'hff) else begin fail = 1; $display("Error 6929: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6930: extop 'h%h !== 1", extop); end
assert (addr === 'hfffef) else begin fail = 1; $display("Error 6931: addr 'h%h !== 'hfffef", addr); end
#2;
clk <= 0;

// f3ffffefffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffefffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1734
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6932: ir 'h%h !== 'hf", ir); end	// Vector No: 1733
assert (op === 'hff) else begin fail = 1; $display("Error 6933: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6934: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6935: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffefffffffff:1:0:b:f8:0:07ffe:
//------------------------

#2;
word <= 'hf3ffffefffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1735
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6936: ir 'h%h !== 'hb", ir); end	// Vector No: 1734
assert (op === 'hf8) else begin fail = 1; $display("Error 6937: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6938: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffe) else begin fail = 1; $display("Error 6939: addr 'h%h !== 'h07ffe", addr); end
#2;
clk <= 0;

// f3ffffefffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffefffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1736
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6940: ir 'h%h !== 'hf", ir); end	// Vector No: 1735
assert (op === 'hf8) else begin fail = 1; $display("Error 6941: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6942: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6943: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffdff3ffffff:0:0:f:ff:0:fffdf:
//------------------------

#2;
word <= 'hffffffdff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1737
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6944: ir 'h%h !== 'hf", ir); end	// Vector No: 1736
assert (op === 'hff) else begin fail = 1; $display("Error 6945: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6946: extop 'h%h !== 0", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 6947: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// ffffffdff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffdff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1738
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6948: ir 'h%h !== 'hf", ir); end	// Vector No: 1737
assert (op === 'hff) else begin fail = 1; $display("Error 6949: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6950: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6951: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffdff3ffffff:1:0:f:f8:0:07ffd:
//------------------------

#2;
word <= 'hffffffdff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1739
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6952: ir 'h%h !== 'hf", ir); end	// Vector No: 1738
assert (op === 'hf8) else begin fail = 1; $display("Error 6953: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6954: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffd) else begin fail = 1; $display("Error 6955: addr 'h%h !== 'h07ffd", addr); end
#2;
clk <= 0;

// ffffffdff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffffdff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1740
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6956: ir 'h%h !== 'hf", ir); end	// Vector No: 1739
assert (op === 'hf0) else begin fail = 1; $display("Error 6957: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6958: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6959: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffdfffffffff:0:0:f:ff:1:fffdf:
//------------------------

#2;
word <= 'hf3ffffdfffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1741
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6960: ir 'h%h !== 'hf", ir); end	// Vector No: 1740
assert (op === 'hff) else begin fail = 1; $display("Error 6961: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6962: extop 'h%h !== 1", extop); end
assert (addr === 'hfffdf) else begin fail = 1; $display("Error 6963: addr 'h%h !== 'hfffdf", addr); end
#2;
clk <= 0;

// f3ffffdfffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffdfffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1742
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6964: ir 'h%h !== 'hf", ir); end	// Vector No: 1741
assert (op === 'hff) else begin fail = 1; $display("Error 6965: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6966: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6967: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffdfffffffff:1:0:b:f8:0:07ffd:
//------------------------

#2;
word <= 'hf3ffffdfffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1743
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 6968: ir 'h%h !== 'hb", ir); end	// Vector No: 1742
assert (op === 'hf8) else begin fail = 1; $display("Error 6969: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6970: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffd) else begin fail = 1; $display("Error 6971: addr 'h%h !== 'h07ffd", addr); end
#2;
clk <= 0;

// f3ffffdfffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffdfffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1744
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6972: ir 'h%h !== 'hf", ir); end	// Vector No: 1743
assert (op === 'hf8) else begin fail = 1; $display("Error 6973: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6974: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 6975: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffffbff3ffffff:0:0:f:ff:0:fffbf:
//------------------------

#2;
word <= 'hffffffbff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1745
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6976: ir 'h%h !== 'hf", ir); end	// Vector No: 1744
assert (op === 'hff) else begin fail = 1; $display("Error 6977: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6978: extop 'h%h !== 0", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 6979: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// ffffffbff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffffbff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1746
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6980: ir 'h%h !== 'hf", ir); end	// Vector No: 1745
assert (op === 'hff) else begin fail = 1; $display("Error 6981: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6982: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6983: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffffbff3ffffff:1:0:f:f8:0:07ffb:
//------------------------

#2;
word <= 'hffffffbff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1747
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6984: ir 'h%h !== 'hf", ir); end	// Vector No: 1746
assert (op === 'hf8) else begin fail = 1; $display("Error 6985: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6986: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffb) else begin fail = 1; $display("Error 6987: addr 'h%h !== 'h07ffb", addr); end
#2;
clk <= 0;

// ffffffbff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffffbff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1748
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6988: ir 'h%h !== 'hf", ir); end	// Vector No: 1747
assert (op === 'hf0) else begin fail = 1; $display("Error 6989: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6990: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 6991: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffbfffffffff:0:0:f:ff:1:fffbf:
//------------------------

#2;
word <= 'hf3ffffbfffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1749
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6992: ir 'h%h !== 'hf", ir); end	// Vector No: 1748
assert (op === 'hff) else begin fail = 1; $display("Error 6993: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 6994: extop 'h%h !== 1", extop); end
assert (addr === 'hfffbf) else begin fail = 1; $display("Error 6995: addr 'h%h !== 'hfffbf", addr); end
#2;
clk <= 0;

// f3ffffbfffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffbfffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1750
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 6996: ir 'h%h !== 'hf", ir); end	// Vector No: 1749
assert (op === 'hff) else begin fail = 1; $display("Error 6997: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 6998: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 6999: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffbfffffffff:1:0:b:f8:0:07ffb:
//------------------------

#2;
word <= 'hf3ffffbfffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1751
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7000: ir 'h%h !== 'hb", ir); end	// Vector No: 1750
assert (op === 'hf8) else begin fail = 1; $display("Error 7001: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7002: extop 'h%h !== 0", extop); end
assert (addr === 'h07ffb) else begin fail = 1; $display("Error 7003: addr 'h%h !== 'h07ffb", addr); end
#2;
clk <= 0;

// f3ffffbfffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffbfffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1752
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7004: ir 'h%h !== 'hf", ir); end	// Vector No: 1751
assert (op === 'hf8) else begin fail = 1; $display("Error 7005: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7006: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7007: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffff7ff3ffffff:0:0:f:ff:0:fff7f:
//------------------------

#2;
word <= 'hffffff7ff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1753
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7008: ir 'h%h !== 'hf", ir); end	// Vector No: 1752
assert (op === 'hff) else begin fail = 1; $display("Error 7009: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7010: extop 'h%h !== 0", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 7011: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// ffffff7ff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffff7ff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1754
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7012: ir 'h%h !== 'hf", ir); end	// Vector No: 1753
assert (op === 'hff) else begin fail = 1; $display("Error 7013: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7014: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7015: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffff7ff3ffffff:1:0:f:f8:0:07ff7:
//------------------------

#2;
word <= 'hffffff7ff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1755
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7016: ir 'h%h !== 'hf", ir); end	// Vector No: 1754
assert (op === 'hf8) else begin fail = 1; $display("Error 7017: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7018: extop 'h%h !== 0", extop); end
assert (addr === 'h07ff7) else begin fail = 1; $display("Error 7019: addr 'h%h !== 'h07ff7", addr); end
#2;
clk <= 0;

// ffffff7ff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffff7ff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1756
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7020: ir 'h%h !== 'hf", ir); end	// Vector No: 1755
assert (op === 'hf0) else begin fail = 1; $display("Error 7021: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7022: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7023: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffff7fffffffff:0:0:f:ff:1:fff7f:
//------------------------

#2;
word <= 'hf3ffff7fffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1757
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7024: ir 'h%h !== 'hf", ir); end	// Vector No: 1756
assert (op === 'hff) else begin fail = 1; $display("Error 7025: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7026: extop 'h%h !== 1", extop); end
assert (addr === 'hfff7f) else begin fail = 1; $display("Error 7027: addr 'h%h !== 'hfff7f", addr); end
#2;
clk <= 0;

// f3ffff7fffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffff7fffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1758
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7028: ir 'h%h !== 'hf", ir); end	// Vector No: 1757
assert (op === 'hff) else begin fail = 1; $display("Error 7029: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7030: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7031: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffff7fffffffff:1:0:b:f8:0:07ff7:
//------------------------

#2;
word <= 'hf3ffff7fffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1759
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7032: ir 'h%h !== 'hb", ir); end	// Vector No: 1758
assert (op === 'hf8) else begin fail = 1; $display("Error 7033: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7034: extop 'h%h !== 0", extop); end
assert (addr === 'h07ff7) else begin fail = 1; $display("Error 7035: addr 'h%h !== 'h07ff7", addr); end
#2;
clk <= 0;

// f3ffff7fffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffff7fffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1760
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7036: ir 'h%h !== 'hf", ir); end	// Vector No: 1759
assert (op === 'hf8) else begin fail = 1; $display("Error 7037: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7038: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7039: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffefff3ffffff:0:0:f:ff:0:ffeff:
//------------------------

#2;
word <= 'hfffffefff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1761
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7040: ir 'h%h !== 'hf", ir); end	// Vector No: 1760
assert (op === 'hff) else begin fail = 1; $display("Error 7041: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7042: extop 'h%h !== 0", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 7043: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// fffffefff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffefff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1762
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7044: ir 'h%h !== 'hf", ir); end	// Vector No: 1761
assert (op === 'hff) else begin fail = 1; $display("Error 7045: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7046: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7047: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffefff3ffffff:1:0:f:f8:0:07fef:
//------------------------

#2;
word <= 'hfffffefff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1763
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7048: ir 'h%h !== 'hf", ir); end	// Vector No: 1762
assert (op === 'hf8) else begin fail = 1; $display("Error 7049: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7050: extop 'h%h !== 0", extop); end
assert (addr === 'h07fef) else begin fail = 1; $display("Error 7051: addr 'h%h !== 'h07fef", addr); end
#2;
clk <= 0;

// fffffefff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffefff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1764
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7052: ir 'h%h !== 'hf", ir); end	// Vector No: 1763
assert (op === 'hf0) else begin fail = 1; $display("Error 7053: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7054: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7055: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffeffffffffff:0:0:f:ff:1:ffeff:
//------------------------

#2;
word <= 'hf3fffeffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1765
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7056: ir 'h%h !== 'hf", ir); end	// Vector No: 1764
assert (op === 'hff) else begin fail = 1; $display("Error 7057: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7058: extop 'h%h !== 1", extop); end
assert (addr === 'hffeff) else begin fail = 1; $display("Error 7059: addr 'h%h !== 'hffeff", addr); end
#2;
clk <= 0;

// f3fffeffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffeffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1766
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7060: ir 'h%h !== 'hf", ir); end	// Vector No: 1765
assert (op === 'hff) else begin fail = 1; $display("Error 7061: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7062: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7063: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffeffffffffff:1:0:b:f8:0:07fef:
//------------------------

#2;
word <= 'hf3fffeffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1767
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7064: ir 'h%h !== 'hb", ir); end	// Vector No: 1766
assert (op === 'hf8) else begin fail = 1; $display("Error 7065: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7066: extop 'h%h !== 0", extop); end
assert (addr === 'h07fef) else begin fail = 1; $display("Error 7067: addr 'h%h !== 'h07fef", addr); end
#2;
clk <= 0;

// f3fffeffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffeffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1768
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7068: ir 'h%h !== 'hf", ir); end	// Vector No: 1767
assert (op === 'hf8) else begin fail = 1; $display("Error 7069: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7070: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7071: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffdfff3ffffff:0:0:f:ff:0:ffdff:
//------------------------

#2;
word <= 'hfffffdfff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1769
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7072: ir 'h%h !== 'hf", ir); end	// Vector No: 1768
assert (op === 'hff) else begin fail = 1; $display("Error 7073: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7074: extop 'h%h !== 0", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 7075: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// fffffdfff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffdfff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1770
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7076: ir 'h%h !== 'hf", ir); end	// Vector No: 1769
assert (op === 'hff) else begin fail = 1; $display("Error 7077: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7078: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7079: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffdfff3ffffff:1:0:f:f8:0:07fdf:
//------------------------

#2;
word <= 'hfffffdfff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1771
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7080: ir 'h%h !== 'hf", ir); end	// Vector No: 1770
assert (op === 'hf8) else begin fail = 1; $display("Error 7081: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7082: extop 'h%h !== 0", extop); end
assert (addr === 'h07fdf) else begin fail = 1; $display("Error 7083: addr 'h%h !== 'h07fdf", addr); end
#2;
clk <= 0;

// fffffdfff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffdfff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1772
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7084: ir 'h%h !== 'hf", ir); end	// Vector No: 1771
assert (op === 'hf0) else begin fail = 1; $display("Error 7085: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7086: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7087: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffdffffffffff:0:0:f:ff:1:ffdff:
//------------------------

#2;
word <= 'hf3fffdffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1773
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7088: ir 'h%h !== 'hf", ir); end	// Vector No: 1772
assert (op === 'hff) else begin fail = 1; $display("Error 7089: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7090: extop 'h%h !== 1", extop); end
assert (addr === 'hffdff) else begin fail = 1; $display("Error 7091: addr 'h%h !== 'hffdff", addr); end
#2;
clk <= 0;

// f3fffdffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffdffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1774
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7092: ir 'h%h !== 'hf", ir); end	// Vector No: 1773
assert (op === 'hff) else begin fail = 1; $display("Error 7093: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7094: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7095: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffdffffffffff:1:0:b:f8:0:07fdf:
//------------------------

#2;
word <= 'hf3fffdffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1775
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7096: ir 'h%h !== 'hb", ir); end	// Vector No: 1774
assert (op === 'hf8) else begin fail = 1; $display("Error 7097: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7098: extop 'h%h !== 0", extop); end
assert (addr === 'h07fdf) else begin fail = 1; $display("Error 7099: addr 'h%h !== 'h07fdf", addr); end
#2;
clk <= 0;

// f3fffdffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffdffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1776
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7100: ir 'h%h !== 'hf", ir); end	// Vector No: 1775
assert (op === 'hf8) else begin fail = 1; $display("Error 7101: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7102: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7103: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffffbfff3ffffff:0:0:f:ff:0:ffbff:
//------------------------

#2;
word <= 'hfffffbfff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1777
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7104: ir 'h%h !== 'hf", ir); end	// Vector No: 1776
assert (op === 'hff) else begin fail = 1; $display("Error 7105: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7106: extop 'h%h !== 0", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 7107: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// fffffbfff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffffbfff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1778
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7108: ir 'h%h !== 'hf", ir); end	// Vector No: 1777
assert (op === 'hff) else begin fail = 1; $display("Error 7109: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7110: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7111: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffffbfff3ffffff:1:0:f:f8:0:07fbf:
//------------------------

#2;
word <= 'hfffffbfff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1779
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7112: ir 'h%h !== 'hf", ir); end	// Vector No: 1778
assert (op === 'hf8) else begin fail = 1; $display("Error 7113: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7114: extop 'h%h !== 0", extop); end
assert (addr === 'h07fbf) else begin fail = 1; $display("Error 7115: addr 'h%h !== 'h07fbf", addr); end
#2;
clk <= 0;

// fffffbfff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffffbfff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1780
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7116: ir 'h%h !== 'hf", ir); end	// Vector No: 1779
assert (op === 'hf0) else begin fail = 1; $display("Error 7117: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7118: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7119: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fffbffffffffff:0:0:f:ff:1:ffbff:
//------------------------

#2;
word <= 'hf3fffbffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1781
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7120: ir 'h%h !== 'hf", ir); end	// Vector No: 1780
assert (op === 'hff) else begin fail = 1; $display("Error 7121: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7122: extop 'h%h !== 1", extop); end
assert (addr === 'hffbff) else begin fail = 1; $display("Error 7123: addr 'h%h !== 'hffbff", addr); end
#2;
clk <= 0;

// f3fffbffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fffbffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1782
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7124: ir 'h%h !== 'hf", ir); end	// Vector No: 1781
assert (op === 'hff) else begin fail = 1; $display("Error 7125: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7126: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7127: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fffbffffffffff:1:0:b:f8:0:07fbf:
//------------------------

#2;
word <= 'hf3fffbffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1783
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7128: ir 'h%h !== 'hb", ir); end	// Vector No: 1782
assert (op === 'hf8) else begin fail = 1; $display("Error 7129: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7130: extop 'h%h !== 0", extop); end
assert (addr === 'h07fbf) else begin fail = 1; $display("Error 7131: addr 'h%h !== 'h07fbf", addr); end
#2;
clk <= 0;

// f3fffbffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fffbffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1784
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7132: ir 'h%h !== 'hf", ir); end	// Vector No: 1783
assert (op === 'hf8) else begin fail = 1; $display("Error 7133: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7134: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7135: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffff7fff3ffffff:0:0:f:ff:0:ff7ff:
//------------------------

#2;
word <= 'hfffff7fff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1785
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7136: ir 'h%h !== 'hf", ir); end	// Vector No: 1784
assert (op === 'hff) else begin fail = 1; $display("Error 7137: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7138: extop 'h%h !== 0", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 7139: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// fffff7fff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffff7fff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1786
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7140: ir 'h%h !== 'hf", ir); end	// Vector No: 1785
assert (op === 'hff) else begin fail = 1; $display("Error 7141: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7142: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7143: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffff7fff3ffffff:1:0:f:f8:0:07f7f:
//------------------------

#2;
word <= 'hfffff7fff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1787
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7144: ir 'h%h !== 'hf", ir); end	// Vector No: 1786
assert (op === 'hf8) else begin fail = 1; $display("Error 7145: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7146: extop 'h%h !== 0", extop); end
assert (addr === 'h07f7f) else begin fail = 1; $display("Error 7147: addr 'h%h !== 'h07f7f", addr); end
#2;
clk <= 0;

// fffff7fff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffff7fff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1788
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7148: ir 'h%h !== 'hf", ir); end	// Vector No: 1787
assert (op === 'hf0) else begin fail = 1; $display("Error 7149: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7150: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7151: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fff7ffffffffff:0:0:f:ff:1:ff7ff:
//------------------------

#2;
word <= 'hf3fff7ffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1789
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7152: ir 'h%h !== 'hf", ir); end	// Vector No: 1788
assert (op === 'hff) else begin fail = 1; $display("Error 7153: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7154: extop 'h%h !== 1", extop); end
assert (addr === 'hff7ff) else begin fail = 1; $display("Error 7155: addr 'h%h !== 'hff7ff", addr); end
#2;
clk <= 0;

// f3fff7ffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fff7ffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1790
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7156: ir 'h%h !== 'hf", ir); end	// Vector No: 1789
assert (op === 'hff) else begin fail = 1; $display("Error 7157: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7158: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7159: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fff7ffffffffff:1:0:b:f8:0:07f7f:
//------------------------

#2;
word <= 'hf3fff7ffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1791
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7160: ir 'h%h !== 'hb", ir); end	// Vector No: 1790
assert (op === 'hf8) else begin fail = 1; $display("Error 7161: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7162: extop 'h%h !== 0", extop); end
assert (addr === 'h07f7f) else begin fail = 1; $display("Error 7163: addr 'h%h !== 'h07f7f", addr); end
#2;
clk <= 0;

// f3fff7ffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fff7ffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1792
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7164: ir 'h%h !== 'hf", ir); end	// Vector No: 1791
assert (op === 'hf8) else begin fail = 1; $display("Error 7165: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7166: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7167: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffeffff3ffffff:0:0:f:ff:0:fefff:
//------------------------

#2;
word <= 'hffffeffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1793
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7168: ir 'h%h !== 'hf", ir); end	// Vector No: 1792
assert (op === 'hff) else begin fail = 1; $display("Error 7169: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7170: extop 'h%h !== 0", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 7171: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// ffffeffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffeffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1794
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7172: ir 'h%h !== 'hf", ir); end	// Vector No: 1793
assert (op === 'hff) else begin fail = 1; $display("Error 7173: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7174: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7175: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffeffff3ffffff:1:0:f:f8:0:07eff:
//------------------------

#2;
word <= 'hffffeffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1795
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7176: ir 'h%h !== 'hf", ir); end	// Vector No: 1794
assert (op === 'hf8) else begin fail = 1; $display("Error 7177: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7178: extop 'h%h !== 0", extop); end
assert (addr === 'h07eff) else begin fail = 1; $display("Error 7179: addr 'h%h !== 'h07eff", addr); end
#2;
clk <= 0;

// ffffeffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffeffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1796
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7180: ir 'h%h !== 'hf", ir); end	// Vector No: 1795
assert (op === 'hf0) else begin fail = 1; $display("Error 7181: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7182: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7183: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffefffffffffff:0:0:f:fe:1:fefff:
//------------------------

#2;
word <= 'hf3ffefffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1797
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7184: ir 'h%h !== 'hf", ir); end	// Vector No: 1796
assert (op === 'hfe) else begin fail = 1; $display("Error 7185: op 'h%h !== 'hfe", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7186: extop 'h%h !== 1", extop); end
assert (addr === 'hfefff) else begin fail = 1; $display("Error 7187: addr 'h%h !== 'hfefff", addr); end
#2;
clk <= 0;

// f3ffefffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffefffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1798
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7188: ir 'h%h !== 'hf", ir); end	// Vector No: 1797
assert (op === 'hff) else begin fail = 1; $display("Error 7189: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7190: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7191: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffefffffffffff:1:0:b:f8:0:07eff:
//------------------------

#2;
word <= 'hf3ffefffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1799
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7192: ir 'h%h !== 'hb", ir); end	// Vector No: 1798
assert (op === 'hf8) else begin fail = 1; $display("Error 7193: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7194: extop 'h%h !== 0", extop); end
assert (addr === 'h07eff) else begin fail = 1; $display("Error 7195: addr 'h%h !== 'h07eff", addr); end
#2;
clk <= 0;

// f3ffefffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffefffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1800
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7196: ir 'h%h !== 'hf", ir); end	// Vector No: 1799
assert (op === 'hf8) else begin fail = 1; $display("Error 7197: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7198: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7199: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffdffff3ffffff:0:0:f:ff:0:fdfff:
//------------------------

#2;
word <= 'hffffdffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1801
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7200: ir 'h%h !== 'hf", ir); end	// Vector No: 1800
assert (op === 'hff) else begin fail = 1; $display("Error 7201: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7202: extop 'h%h !== 0", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 7203: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// ffffdffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffdffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1802
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7204: ir 'h%h !== 'hf", ir); end	// Vector No: 1801
assert (op === 'hff) else begin fail = 1; $display("Error 7205: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7206: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7207: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffdffff3ffffff:1:0:f:f8:0:07dff:
//------------------------

#2;
word <= 'hffffdffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1803
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7208: ir 'h%h !== 'hf", ir); end	// Vector No: 1802
assert (op === 'hf8) else begin fail = 1; $display("Error 7209: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7210: extop 'h%h !== 0", extop); end
assert (addr === 'h07dff) else begin fail = 1; $display("Error 7211: addr 'h%h !== 'h07dff", addr); end
#2;
clk <= 0;

// ffffdffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffdffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1804
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7212: ir 'h%h !== 'hf", ir); end	// Vector No: 1803
assert (op === 'hf0) else begin fail = 1; $display("Error 7213: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7214: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7215: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffdfffffffffff:0:0:f:fd:1:fdfff:
//------------------------

#2;
word <= 'hf3ffdfffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1805
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7216: ir 'h%h !== 'hf", ir); end	// Vector No: 1804
assert (op === 'hfd) else begin fail = 1; $display("Error 7217: op 'h%h !== 'hfd", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7218: extop 'h%h !== 1", extop); end
assert (addr === 'hfdfff) else begin fail = 1; $display("Error 7219: addr 'h%h !== 'hfdfff", addr); end
#2;
clk <= 0;

// f3ffdfffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffdfffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1806
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7220: ir 'h%h !== 'hf", ir); end	// Vector No: 1805
assert (op === 'hff) else begin fail = 1; $display("Error 7221: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7222: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7223: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffdfffffffffff:1:0:b:f8:0:07dff:
//------------------------

#2;
word <= 'hf3ffdfffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1807
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7224: ir 'h%h !== 'hb", ir); end	// Vector No: 1806
assert (op === 'hf8) else begin fail = 1; $display("Error 7225: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7226: extop 'h%h !== 0", extop); end
assert (addr === 'h07dff) else begin fail = 1; $display("Error 7227: addr 'h%h !== 'h07dff", addr); end
#2;
clk <= 0;

// f3ffdfffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffdfffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1808
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7228: ir 'h%h !== 'hf", ir); end	// Vector No: 1807
assert (op === 'hf8) else begin fail = 1; $display("Error 7229: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7230: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7231: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffffbffff3ffffff:0:0:f:ff:0:fbfff:
//------------------------

#2;
word <= 'hffffbffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1809
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7232: ir 'h%h !== 'hf", ir); end	// Vector No: 1808
assert (op === 'hff) else begin fail = 1; $display("Error 7233: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7234: extop 'h%h !== 0", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 7235: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// ffffbffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffffbffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1810
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7236: ir 'h%h !== 'hf", ir); end	// Vector No: 1809
assert (op === 'hff) else begin fail = 1; $display("Error 7237: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7238: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7239: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffffbffff3ffffff:1:0:f:f8:0:07bff:
//------------------------

#2;
word <= 'hffffbffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1811
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7240: ir 'h%h !== 'hf", ir); end	// Vector No: 1810
assert (op === 'hf8) else begin fail = 1; $display("Error 7241: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7242: extop 'h%h !== 0", extop); end
assert (addr === 'h07bff) else begin fail = 1; $display("Error 7243: addr 'h%h !== 'h07bff", addr); end
#2;
clk <= 0;

// ffffbffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffffbffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1812
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7244: ir 'h%h !== 'hf", ir); end	// Vector No: 1811
assert (op === 'hf0) else begin fail = 1; $display("Error 7245: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7246: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7247: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffbfffffffffff:0:0:f:fb:1:fbfff:
//------------------------

#2;
word <= 'hf3ffbfffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1813
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7248: ir 'h%h !== 'hf", ir); end	// Vector No: 1812
assert (op === 'hfb) else begin fail = 1; $display("Error 7249: op 'h%h !== 'hfb", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7250: extop 'h%h !== 1", extop); end
assert (addr === 'hfbfff) else begin fail = 1; $display("Error 7251: addr 'h%h !== 'hfbfff", addr); end
#2;
clk <= 0;

// f3ffbfffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffbfffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1814
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7252: ir 'h%h !== 'hf", ir); end	// Vector No: 1813
assert (op === 'hff) else begin fail = 1; $display("Error 7253: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7254: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7255: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffbfffffffffff:1:0:b:f8:0:07bff:
//------------------------

#2;
word <= 'hf3ffbfffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1815
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7256: ir 'h%h !== 'hb", ir); end	// Vector No: 1814
assert (op === 'hf8) else begin fail = 1; $display("Error 7257: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7258: extop 'h%h !== 0", extop); end
assert (addr === 'h07bff) else begin fail = 1; $display("Error 7259: addr 'h%h !== 'h07bff", addr); end
#2;
clk <= 0;

// f3ffbfffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffbfffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1816
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7260: ir 'h%h !== 'hf", ir); end	// Vector No: 1815
assert (op === 'hf8) else begin fail = 1; $display("Error 7261: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7262: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7263: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffff7ffff3ffffff:0:0:f:ff:0:f7fff:
//------------------------

#2;
word <= 'hffff7ffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1817
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7264: ir 'h%h !== 'hf", ir); end	// Vector No: 1816
assert (op === 'hff) else begin fail = 1; $display("Error 7265: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7266: extop 'h%h !== 0", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 7267: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// ffff7ffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffff7ffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1818
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7268: ir 'h%h !== 'hf", ir); end	// Vector No: 1817
assert (op === 'hff) else begin fail = 1; $display("Error 7269: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7270: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7271: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffff7ffff3ffffff:1:0:f:f8:0:077ff:
//------------------------

#2;
word <= 'hffff7ffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1819
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7272: ir 'h%h !== 'hf", ir); end	// Vector No: 1818
assert (op === 'hf8) else begin fail = 1; $display("Error 7273: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7274: extop 'h%h !== 0", extop); end
assert (addr === 'h077ff) else begin fail = 1; $display("Error 7275: addr 'h%h !== 'h077ff", addr); end
#2;
clk <= 0;

// ffff7ffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffff7ffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1820
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7276: ir 'h%h !== 'hf", ir); end	// Vector No: 1819
assert (op === 'hf0) else begin fail = 1; $display("Error 7277: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7278: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7279: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ff7fffffffffff:0:0:f:f7:1:f7fff:
//------------------------

#2;
word <= 'hf3ff7fffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1821
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7280: ir 'h%h !== 'hf", ir); end	// Vector No: 1820
assert (op === 'hf7) else begin fail = 1; $display("Error 7281: op 'h%h !== 'hf7", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7282: extop 'h%h !== 1", extop); end
assert (addr === 'hf7fff) else begin fail = 1; $display("Error 7283: addr 'h%h !== 'hf7fff", addr); end
#2;
clk <= 0;

// f3ff7fffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ff7fffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1822
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7284: ir 'h%h !== 'hf", ir); end	// Vector No: 1821
assert (op === 'hff) else begin fail = 1; $display("Error 7285: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7286: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7287: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ff7fffffffffff:1:0:b:f8:0:077ff:
//------------------------

#2;
word <= 'hf3ff7fffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1823
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7288: ir 'h%h !== 'hb", ir); end	// Vector No: 1822
assert (op === 'hf8) else begin fail = 1; $display("Error 7289: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7290: extop 'h%h !== 0", extop); end
assert (addr === 'h077ff) else begin fail = 1; $display("Error 7291: addr 'h%h !== 'h077ff", addr); end
#2;
clk <= 0;

// f3ff7fffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ff7fffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1824
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7292: ir 'h%h !== 'hf", ir); end	// Vector No: 1823
assert (op === 'hf8) else begin fail = 1; $display("Error 7293: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7294: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7295: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffefffff3ffffff:0:0:f:ff:0:effff:
//------------------------

#2;
word <= 'hfffefffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1825
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7296: ir 'h%h !== 'hf", ir); end	// Vector No: 1824
assert (op === 'hff) else begin fail = 1; $display("Error 7297: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7298: extop 'h%h !== 0", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 7299: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// fffefffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffefffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1826
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7300: ir 'h%h !== 'hf", ir); end	// Vector No: 1825
assert (op === 'hff) else begin fail = 1; $display("Error 7301: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7302: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7303: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffefffff3ffffff:1:0:f:f8:0:06fff:
//------------------------

#2;
word <= 'hfffefffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1827
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7304: ir 'h%h !== 'hf", ir); end	// Vector No: 1826
assert (op === 'hf8) else begin fail = 1; $display("Error 7305: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7306: extop 'h%h !== 0", extop); end
assert (addr === 'h06fff) else begin fail = 1; $display("Error 7307: addr 'h%h !== 'h06fff", addr); end
#2;
clk <= 0;

// fffefffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffefffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1828
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7308: ir 'h%h !== 'hf", ir); end	// Vector No: 1827
assert (op === 'hf0) else begin fail = 1; $display("Error 7309: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7310: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7311: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3feffffffffffff:0:0:f:ef:1:effff:
//------------------------

#2;
word <= 'hf3feffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1829
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7312: ir 'h%h !== 'hf", ir); end	// Vector No: 1828
assert (op === 'hef) else begin fail = 1; $display("Error 7313: op 'h%h !== 'hef", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7314: extop 'h%h !== 1", extop); end
assert (addr === 'heffff) else begin fail = 1; $display("Error 7315: addr 'h%h !== 'heffff", addr); end
#2;
clk <= 0;

// f3feffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3feffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1830
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7316: ir 'h%h !== 'hf", ir); end	// Vector No: 1829
assert (op === 'hff) else begin fail = 1; $display("Error 7317: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7318: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7319: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3feffffffffffff:1:0:b:f8:0:06fff:
//------------------------

#2;
word <= 'hf3feffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1831
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7320: ir 'h%h !== 'hb", ir); end	// Vector No: 1830
assert (op === 'hf8) else begin fail = 1; $display("Error 7321: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7322: extop 'h%h !== 0", extop); end
assert (addr === 'h06fff) else begin fail = 1; $display("Error 7323: addr 'h%h !== 'h06fff", addr); end
#2;
clk <= 0;

// f3feffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3feffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1832
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7324: ir 'h%h !== 'hf", ir); end	// Vector No: 1831
assert (op === 'hf8) else begin fail = 1; $display("Error 7325: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7326: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7327: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffdfffff3ffffff:0:0:f:ff:0:dffff:
//------------------------

#2;
word <= 'hfffdfffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1833
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7328: ir 'h%h !== 'hf", ir); end	// Vector No: 1832
assert (op === 'hff) else begin fail = 1; $display("Error 7329: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7330: extop 'h%h !== 0", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 7331: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// fffdfffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffdfffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1834
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7332: ir 'h%h !== 'hf", ir); end	// Vector No: 1833
assert (op === 'hff) else begin fail = 1; $display("Error 7333: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7334: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7335: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffdfffff3ffffff:1:0:f:f8:0:05fff:
//------------------------

#2;
word <= 'hfffdfffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1835
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7336: ir 'h%h !== 'hf", ir); end	// Vector No: 1834
assert (op === 'hf8) else begin fail = 1; $display("Error 7337: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7338: extop 'h%h !== 0", extop); end
assert (addr === 'h05fff) else begin fail = 1; $display("Error 7339: addr 'h%h !== 'h05fff", addr); end
#2;
clk <= 0;

// fffdfffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffdfffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1836
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7340: ir 'h%h !== 'hf", ir); end	// Vector No: 1835
assert (op === 'hf0) else begin fail = 1; $display("Error 7341: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7342: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7343: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fdffffffffffff:0:0:f:df:1:dffff:
//------------------------

#2;
word <= 'hf3fdffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1837
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7344: ir 'h%h !== 'hf", ir); end	// Vector No: 1836
assert (op === 'hdf) else begin fail = 1; $display("Error 7345: op 'h%h !== 'hdf", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7346: extop 'h%h !== 1", extop); end
assert (addr === 'hdffff) else begin fail = 1; $display("Error 7347: addr 'h%h !== 'hdffff", addr); end
#2;
clk <= 0;

// f3fdffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fdffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1838
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7348: ir 'h%h !== 'hf", ir); end	// Vector No: 1837
assert (op === 'hff) else begin fail = 1; $display("Error 7349: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7350: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7351: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fdffffffffffff:1:0:b:f8:0:05fff:
//------------------------

#2;
word <= 'hf3fdffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1839
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7352: ir 'h%h !== 'hb", ir); end	// Vector No: 1838
assert (op === 'hf8) else begin fail = 1; $display("Error 7353: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7354: extop 'h%h !== 0", extop); end
assert (addr === 'h05fff) else begin fail = 1; $display("Error 7355: addr 'h%h !== 'h05fff", addr); end
#2;
clk <= 0;

// f3fdffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fdffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1840
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7356: ir 'h%h !== 'hf", ir); end	// Vector No: 1839
assert (op === 'hf8) else begin fail = 1; $display("Error 7357: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7358: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7359: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fffbfffff3ffffff:0:0:f:ff:0:bffff:
//------------------------

#2;
word <= 'hfffbfffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1841
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7360: ir 'h%h !== 'hf", ir); end	// Vector No: 1840
assert (op === 'hff) else begin fail = 1; $display("Error 7361: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7362: extop 'h%h !== 0", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 7363: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// fffbfffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfffbfffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1842
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7364: ir 'h%h !== 'hf", ir); end	// Vector No: 1841
assert (op === 'hff) else begin fail = 1; $display("Error 7365: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7366: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7367: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fffbfffff3ffffff:1:0:f:f8:0:03fff:
//------------------------

#2;
word <= 'hfffbfffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1843
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7368: ir 'h%h !== 'hf", ir); end	// Vector No: 1842
assert (op === 'hf8) else begin fail = 1; $display("Error 7369: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7370: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7371: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fffbfffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfffbfffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1844
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7372: ir 'h%h !== 'hf", ir); end	// Vector No: 1843
assert (op === 'hf0) else begin fail = 1; $display("Error 7373: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7374: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7375: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fbffffffffffff:0:0:f:bf:1:bffff:
//------------------------

#2;
word <= 'hf3fbffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1845
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7376: ir 'h%h !== 'hf", ir); end	// Vector No: 1844
assert (op === 'hbf) else begin fail = 1; $display("Error 7377: op 'h%h !== 'hbf", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7378: extop 'h%h !== 1", extop); end
assert (addr === 'hbffff) else begin fail = 1; $display("Error 7379: addr 'h%h !== 'hbffff", addr); end
#2;
clk <= 0;

// f3fbffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3fbffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1846
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7380: ir 'h%h !== 'hf", ir); end	// Vector No: 1845
assert (op === 'hff) else begin fail = 1; $display("Error 7381: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7382: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7383: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3fbffffffffffff:1:0:b:f8:0:03fff:
//------------------------

#2;
word <= 'hf3fbffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1847
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7384: ir 'h%h !== 'hb", ir); end	// Vector No: 1846
assert (op === 'hf8) else begin fail = 1; $display("Error 7385: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7386: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7387: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3fbffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3fbffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1848
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7388: ir 'h%h !== 'hf", ir); end	// Vector No: 1847
assert (op === 'hf8) else begin fail = 1; $display("Error 7389: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7390: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7391: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fff7fffff3ffffff:0:0:f:ff:0:7ffff:
//------------------------

#2;
word <= 'hfff7fffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1849
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7392: ir 'h%h !== 'hf", ir); end	// Vector No: 1848
assert (op === 'hff) else begin fail = 1; $display("Error 7393: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7394: extop 'h%h !== 0", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 7395: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// fff7fffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfff7fffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1850
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7396: ir 'h%h !== 'hf", ir); end	// Vector No: 1849
assert (op === 'hff) else begin fail = 1; $display("Error 7397: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7398: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7399: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fff7fffff3ffffff:1:0:f:f0:0:07fff:
//------------------------

#2;
word <= 'hfff7fffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1851
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7400: ir 'h%h !== 'hf", ir); end	// Vector No: 1850
assert (op === 'hf0) else begin fail = 1; $display("Error 7401: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7402: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7403: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fff7fffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfff7fffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1852
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7404: ir 'h%h !== 'hf", ir); end	// Vector No: 1851
assert (op === 'hf0) else begin fail = 1; $display("Error 7405: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7406: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7407: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3f7ffffffffffff:0:0:f:7f:1:7ffff:
//------------------------

#2;
word <= 'hf3f7ffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1853
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7408: ir 'h%h !== 'hf", ir); end	// Vector No: 1852
assert (op === 'h7f) else begin fail = 1; $display("Error 7409: op 'h%h !== 'h7f", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7410: extop 'h%h !== 1", extop); end
assert (addr === 'h7ffff) else begin fail = 1; $display("Error 7411: addr 'h%h !== 'h7ffff", addr); end
#2;
clk <= 0;

// f3f7ffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3f7ffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1854
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7412: ir 'h%h !== 'hf", ir); end	// Vector No: 1853
assert (op === 'hff) else begin fail = 1; $display("Error 7413: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7414: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7415: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3f7ffffffffffff:1:0:b:f0:0:07fff:
//------------------------

#2;
word <= 'hf3f7ffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1855
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7416: ir 'h%h !== 'hb", ir); end	// Vector No: 1854
assert (op === 'hf0) else begin fail = 1; $display("Error 7417: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7418: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7419: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3f7ffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3f7ffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1856
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7420: ir 'h%h !== 'hf", ir); end	// Vector No: 1855
assert (op === 'hf8) else begin fail = 1; $display("Error 7421: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7422: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7423: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffeffffff3ffffff:0:0:f:fe:0:fffff:
//------------------------

#2;
word <= 'hffeffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1857
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7424: ir 'h%h !== 'hf", ir); end	// Vector No: 1856
assert (op === 'hfe) else begin fail = 1; $display("Error 7425: op 'h%h !== 'hfe", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7426: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7427: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffeffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffeffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1858
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7428: ir 'h%h !== 'hf", ir); end	// Vector No: 1857
assert (op === 'hff) else begin fail = 1; $display("Error 7429: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7430: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7431: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffeffffff3ffffff:1:0:f:e8:0:07fff:
//------------------------

#2;
word <= 'hffeffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1859
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7432: ir 'h%h !== 'hf", ir); end	// Vector No: 1858
assert (op === 'he8) else begin fail = 1; $display("Error 7433: op 'h%h !== 'he8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7434: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7435: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffeffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffeffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1860
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7436: ir 'h%h !== 'hf", ir); end	// Vector No: 1859
assert (op === 'hf0) else begin fail = 1; $display("Error 7437: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7438: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7439: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffff:0:0:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1861
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7440: ir 'h%h !== 'hf", ir); end	// Vector No: 1860
assert (op === 'hff) else begin fail = 1; $display("Error 7441: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7442: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7443: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hf3ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1862
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7444: ir 'h%h !== 'hf", ir); end	// Vector No: 1861
assert (op === 'hff) else begin fail = 1; $display("Error 7445: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7446: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7447: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f3ffffffffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1863
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7448: ir 'h%h !== 'hb", ir); end	// Vector No: 1862
assert (op === 'hf8) else begin fail = 1; $display("Error 7449: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7450: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7451: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f3ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf3ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1864
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7452: ir 'h%h !== 'hf", ir); end	// Vector No: 1863
assert (op === 'hf8) else begin fail = 1; $display("Error 7453: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7454: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7455: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffdffffff3ffffff:0:0:f:fd:0:fffff:
//------------------------

#2;
word <= 'hffdffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1865
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7456: ir 'h%h !== 'hf", ir); end	// Vector No: 1864
assert (op === 'hfd) else begin fail = 1; $display("Error 7457: op 'h%h !== 'hfd", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7458: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7459: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffdffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffdffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1866
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7460: ir 'h%h !== 'hf", ir); end	// Vector No: 1865
assert (op === 'hff) else begin fail = 1; $display("Error 7461: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7462: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7463: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffdffffff3ffffff:1:0:f:d8:0:07fff:
//------------------------

#2;
word <= 'hffdffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1867
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7464: ir 'h%h !== 'hf", ir); end	// Vector No: 1866
assert (op === 'hd8) else begin fail = 1; $display("Error 7465: op 'h%h !== 'hd8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7466: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7467: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffdffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffdffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1868
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7468: ir 'h%h !== 'hf", ir); end	// Vector No: 1867
assert (op === 'hf0) else begin fail = 1; $display("Error 7469: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7470: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7471: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// ffbffffff3ffffff:0:0:f:fb:0:fffff:
//------------------------

#2;
word <= 'hffbffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1869
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7472: ir 'h%h !== 'hf", ir); end	// Vector No: 1868
assert (op === 'hfb) else begin fail = 1; $display("Error 7473: op 'h%h !== 'hfb", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7474: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7475: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffbffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hffbffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1870
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7476: ir 'h%h !== 'hf", ir); end	// Vector No: 1869
assert (op === 'hff) else begin fail = 1; $display("Error 7477: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7478: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7479: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ffbffffff3ffffff:1:0:f:b8:0:07fff:
//------------------------

#2;
word <= 'hffbffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1871
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7480: ir 'h%h !== 'hf", ir); end	// Vector No: 1870
assert (op === 'hb8) else begin fail = 1; $display("Error 7481: op 'h%h !== 'hb8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7482: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7483: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ffbffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hffbffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1872
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7484: ir 'h%h !== 'hf", ir); end	// Vector No: 1871
assert (op === 'hf0) else begin fail = 1; $display("Error 7485: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7486: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7487: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// ff7ffffff3ffffff:0:0:f:f7:0:fffff:
//------------------------

#2;
word <= 'hff7ffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1873
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7488: ir 'h%h !== 'hf", ir); end	// Vector No: 1872
assert (op === 'hf7) else begin fail = 1; $display("Error 7489: op 'h%h !== 'hf7", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7490: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7491: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ff7ffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hff7ffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1874
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7492: ir 'h%h !== 'hf", ir); end	// Vector No: 1873
assert (op === 'hff) else begin fail = 1; $display("Error 7493: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7494: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7495: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// ff7ffffff3ffffff:1:0:f:7f:0:07fff:
//------------------------

#2;
word <= 'hff7ffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1875
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7496: ir 'h%h !== 'hf", ir); end	// Vector No: 1874
assert (op === 'h7f) else begin fail = 1; $display("Error 7497: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7498: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7499: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// ff7ffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hff7ffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1876
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7500: ir 'h%h !== 'hf", ir); end	// Vector No: 1875
assert (op === 'hf0) else begin fail = 1; $display("Error 7501: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7502: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7503: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fefffffff3ffffff:0:0:f:ef:0:fffff:
//------------------------

#2;
word <= 'hfefffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1877
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7504: ir 'h%h !== 'hf", ir); end	// Vector No: 1876
assert (op === 'hef) else begin fail = 1; $display("Error 7505: op 'h%h !== 'hef", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7506: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7507: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fefffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfefffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1878
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7508: ir 'h%h !== 'hf", ir); end	// Vector No: 1877
assert (op === 'hff) else begin fail = 1; $display("Error 7509: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7510: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7511: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fefffffff3ffffff:1:0:e:f8:0:07fff:
//------------------------

#2;
word <= 'hfefffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1879
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 7512: ir 'h%h !== 'he", ir); end	// Vector No: 1878
assert (op === 'hf8) else begin fail = 1; $display("Error 7513: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7514: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7515: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fefffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfefffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1880
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7516: ir 'h%h !== 'hf", ir); end	// Vector No: 1879
assert (op === 'hf0) else begin fail = 1; $display("Error 7517: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7518: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7519: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fdfffffff3ffffff:0:0:f:df:0:fffff:
//------------------------

#2;
word <= 'hfdfffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1881
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7520: ir 'h%h !== 'hf", ir); end	// Vector No: 1880
assert (op === 'hdf) else begin fail = 1; $display("Error 7521: op 'h%h !== 'hdf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7522: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7523: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fdfffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfdfffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1882
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7524: ir 'h%h !== 'hf", ir); end	// Vector No: 1881
assert (op === 'hff) else begin fail = 1; $display("Error 7525: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7526: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7527: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fdfffffff3ffffff:1:0:d:f8:0:07fff:
//------------------------

#2;
word <= 'hfdfffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1883
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 7528: ir 'h%h !== 'hd", ir); end	// Vector No: 1882
assert (op === 'hf8) else begin fail = 1; $display("Error 7529: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7530: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7531: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fdfffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfdfffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1884
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7532: ir 'h%h !== 'hf", ir); end	// Vector No: 1883
assert (op === 'hf0) else begin fail = 1; $display("Error 7533: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7534: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7535: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// fbfffffff3ffffff:0:0:f:bf:0:fffff:
//------------------------

#2;
word <= 'hfbfffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1885
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7536: ir 'h%h !== 'hf", ir); end	// Vector No: 1884
assert (op === 'hbf) else begin fail = 1; $display("Error 7537: op 'h%h !== 'hbf", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7538: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7539: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fbfffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hfbfffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1886
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7540: ir 'h%h !== 'hf", ir); end	// Vector No: 1885
assert (op === 'hff) else begin fail = 1; $display("Error 7541: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7542: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7543: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// fbfffffff3ffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hfbfffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1887
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7544: ir 'h%h !== 'hb", ir); end	// Vector No: 1886
assert (op === 'hf8) else begin fail = 1; $display("Error 7545: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7546: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7547: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// fbfffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hfbfffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1888
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7548: ir 'h%h !== 'hf", ir); end	// Vector No: 1887
assert (op === 'hf0) else begin fail = 1; $display("Error 7549: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7550: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7551: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// f7fffffff3ffffff:0:0:f:7f:0:fffff:
//------------------------

#2;
word <= 'hf7fffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1889
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7552: ir 'h%h !== 'hf", ir); end	// Vector No: 1888
assert (op === 'h7f) else begin fail = 1; $display("Error 7553: op 'h%h !== 'h7f", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7554: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7555: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f7fffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hf7fffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1890
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7556: ir 'h%h !== 'hf", ir); end	// Vector No: 1889
assert (op === 'hff) else begin fail = 1; $display("Error 7557: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7558: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7559: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// f7fffffff3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hf7fffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1891
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7560: ir 'h%h !== 'hf", ir); end	// Vector No: 1890
assert (op === 'hf8) else begin fail = 1; $display("Error 7561: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7562: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7563: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// f7fffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hf7fffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1892
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7564: ir 'h%h !== 'hf", ir); end	// Vector No: 1891
assert (op === 'hf0) else begin fail = 1; $display("Error 7565: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7566: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7567: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// effffffff3ffffff:0:0:e:ff:0:fffff:
//------------------------

#2;
word <= 'heffffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1893
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 7568: ir 'h%h !== 'he", ir); end	// Vector No: 1892
assert (op === 'hff) else begin fail = 1; $display("Error 7569: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7570: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7571: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// effffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'heffffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1894
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7572: ir 'h%h !== 'hf", ir); end	// Vector No: 1893
assert (op === 'hff) else begin fail = 1; $display("Error 7573: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7574: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7575: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// effffffff3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'heffffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1895
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7576: ir 'h%h !== 'hf", ir); end	// Vector No: 1894
assert (op === 'hf8) else begin fail = 1; $display("Error 7577: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7578: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7579: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// effffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'heffffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1896
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7580: ir 'h%h !== 'hf", ir); end	// Vector No: 1895
assert (op === 'hf0) else begin fail = 1; $display("Error 7581: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7582: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7583: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// e3ffffffffffffff:0:0:e:ff:1:fffff:
//------------------------

#2;
word <= 'he3ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1897
#2;

assert (ir === 'he) else begin fail = 1; $display("Error 7584: ir 'h%h !== 'he", ir); end	// Vector No: 1896
assert (op === 'hff) else begin fail = 1; $display("Error 7585: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7586: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7587: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// e3ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'he3ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1898
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7588: ir 'h%h !== 'hf", ir); end	// Vector No: 1897
assert (op === 'hff) else begin fail = 1; $display("Error 7589: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7590: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7591: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// e3ffffffffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'he3ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1899
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7592: ir 'h%h !== 'hb", ir); end	// Vector No: 1898
assert (op === 'hf8) else begin fail = 1; $display("Error 7593: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7594: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7595: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// e3ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'he3ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1900
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7596: ir 'h%h !== 'hf", ir); end	// Vector No: 1899
assert (op === 'hf8) else begin fail = 1; $display("Error 7597: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7598: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7599: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// dffffffff3ffffff:0:0:d:ff:0:fffff:
//------------------------

#2;
word <= 'hdffffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1901
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 7600: ir 'h%h !== 'hd", ir); end	// Vector No: 1900
assert (op === 'hff) else begin fail = 1; $display("Error 7601: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7602: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7603: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// dffffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hdffffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1902
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7604: ir 'h%h !== 'hf", ir); end	// Vector No: 1901
assert (op === 'hff) else begin fail = 1; $display("Error 7605: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7606: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7607: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// dffffffff3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hdffffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1903
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7608: ir 'h%h !== 'hf", ir); end	// Vector No: 1902
assert (op === 'hf8) else begin fail = 1; $display("Error 7609: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7610: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7611: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// dffffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hdffffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1904
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7612: ir 'h%h !== 'hf", ir); end	// Vector No: 1903
assert (op === 'hf0) else begin fail = 1; $display("Error 7613: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7614: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7615: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// d3ffffffffffffff:0:0:d:ff:1:fffff:
//------------------------

#2;
word <= 'hd3ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1905
#2;

assert (ir === 'hd) else begin fail = 1; $display("Error 7616: ir 'h%h !== 'hd", ir); end	// Vector No: 1904
assert (op === 'hff) else begin fail = 1; $display("Error 7617: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7618: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7619: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// d3ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hd3ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1906
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7620: ir 'h%h !== 'hf", ir); end	// Vector No: 1905
assert (op === 'hff) else begin fail = 1; $display("Error 7621: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7622: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7623: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// d3ffffffffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hd3ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1907
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7624: ir 'h%h !== 'hb", ir); end	// Vector No: 1906
assert (op === 'hf8) else begin fail = 1; $display("Error 7625: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7626: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7627: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// d3ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hd3ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1908
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7628: ir 'h%h !== 'hf", ir); end	// Vector No: 1907
assert (op === 'hf8) else begin fail = 1; $display("Error 7629: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7630: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7631: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// bffffffff3ffffff:0:0:b:ff:0:fffff:
//------------------------

#2;
word <= 'hbffffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1909
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7632: ir 'h%h !== 'hb", ir); end	// Vector No: 1908
assert (op === 'hff) else begin fail = 1; $display("Error 7633: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7634: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7635: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// bffffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'hbffffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1910
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7636: ir 'h%h !== 'hf", ir); end	// Vector No: 1909
assert (op === 'hff) else begin fail = 1; $display("Error 7637: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7638: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7639: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// bffffffff3ffffff:1:0:f:f8:0:07fff:
//------------------------

#2;
word <= 'hbffffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1911
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7640: ir 'h%h !== 'hf", ir); end	// Vector No: 1910
assert (op === 'hf8) else begin fail = 1; $display("Error 7641: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7642: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7643: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// bffffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'hbffffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1912
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7644: ir 'h%h !== 'hf", ir); end	// Vector No: 1911
assert (op === 'hf0) else begin fail = 1; $display("Error 7645: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7646: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7647: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// b3ffffffffffffff:0:0:b:ff:1:fffff:
//------------------------

#2;
word <= 'hb3ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1913
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7648: ir 'h%h !== 'hb", ir); end	// Vector No: 1912
assert (op === 'hff) else begin fail = 1; $display("Error 7649: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7650: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7651: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// b3ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'hb3ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1914
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7652: ir 'h%h !== 'hf", ir); end	// Vector No: 1913
assert (op === 'hff) else begin fail = 1; $display("Error 7653: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7654: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7655: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// b3ffffffffffffff:1:0:b:f8:0:07fff:
//------------------------

#2;
word <= 'hb3ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1915
#2;

assert (ir === 'hb) else begin fail = 1; $display("Error 7656: ir 'h%h !== 'hb", ir); end	// Vector No: 1914
assert (op === 'hf8) else begin fail = 1; $display("Error 7657: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7658: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7659: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// b3ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'hb3ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1916
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7660: ir 'h%h !== 'hf", ir); end	// Vector No: 1915
assert (op === 'hf8) else begin fail = 1; $display("Error 7661: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7662: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7663: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 7ffffffff3ffffff:0:0:7:ff:0:fffff:
//------------------------

#2;
word <= 'h7ffffffff3ffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1917
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 7664: ir 'h%h !== 'h7", ir); end	// Vector No: 1916
assert (op === 'hff) else begin fail = 1; $display("Error 7665: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7666: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7667: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 7ffffffff3ffffff:0:1:f:ff:1:fffff:
//------------------------

#2;
word <= 'h7ffffffff3ffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1918
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7668: ir 'h%h !== 'hf", ir); end	// Vector No: 1917
assert (op === 'hff) else begin fail = 1; $display("Error 7669: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7670: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7671: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 7ffffffff3ffffff:1:0:7:f8:0:07fff:
//------------------------

#2;
word <= 'h7ffffffff3ffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1919
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 7672: ir 'h%h !== 'h7", ir); end	// Vector No: 1918
assert (op === 'hf8) else begin fail = 1; $display("Error 7673: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7674: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7675: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 7ffffffff3ffffff:1:1:f:f0:0:03fff:
//------------------------

#2;
word <= 'h7ffffffff3ffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1920
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7676: ir 'h%h !== 'hf", ir); end	// Vector No: 1919
assert (op === 'hf0) else begin fail = 1; $display("Error 7677: op 'h%h !== 'hf0", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7678: extop 'h%h !== 0", extop); end
assert (addr === 'h03fff) else begin fail = 1; $display("Error 7679: addr 'h%h !== 'h03fff", addr); end
#2;
clk <= 0;

// 73ffffffffffffff:0:0:7:ff:1:fffff:
//------------------------

#2;
word <= 'h73ffffffffffffff;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1921
#2;

assert (ir === 'h7) else begin fail = 1; $display("Error 7680: ir 'h%h !== 'h7", ir); end	// Vector No: 1920
assert (op === 'hff) else begin fail = 1; $display("Error 7681: op 'h%h !== 'hff", op); end
assert (extop === 1) else begin fail = 1; $display("Error 7682: extop 'h%h !== 1", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7683: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 73ffffffffffffff:0:1:f:ff:0:fffff:
//------------------------

#2;
word <= 'h73ffffffffffffff;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1922
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7684: ir 'h%h !== 'hf", ir); end	// Vector No: 1921
assert (op === 'hff) else begin fail = 1; $display("Error 7685: op 'h%h !== 'hff", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7686: extop 'h%h !== 0", extop); end
assert (addr === 'hfffff) else begin fail = 1; $display("Error 7687: addr 'h%h !== 'hfffff", addr); end
#2;
clk <= 0;

// 73ffffffffffffff:1:0:3:f8:0:07fff:
//------------------------

#2;
word <= 'h73ffffffffffffff;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1923
#2;

assert (ir === 'h3) else begin fail = 1; $display("Error 7688: ir 'h%h !== 'h3", ir); end	// Vector No: 1922
assert (op === 'hf8) else begin fail = 1; $display("Error 7689: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7690: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7691: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

// 73ffffffffffffff:1:1:f:f8:0:07fff:
//------------------------

#2;
word <= 'h73ffffffffffffff;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1924
#2;

assert (ir === 'hf) else begin fail = 1; $display("Error 7692: ir 'h%h !== 'hf", ir); end	// Vector No: 1923
assert (op === 'hf8) else begin fail = 1; $display("Error 7693: op 'h%h !== 'hf8", op); end
assert (extop === 0) else begin fail = 1; $display("Error 7694: extop 'h%h !== 0", extop); end
assert (addr === 'h07fff) else begin fail = 1; $display("Error 7695: addr 'h%h !== 'h07fff", addr); end
#2;
clk <= 0;

#4;
if (fail) begin
    $display("Test FAIL");
    $display("------------------------");
    $finish(1);
end
$display("Test PASS");
$display("------------------------");
$finish;

end

endmodule
