// ALU:
// ALUS -> I[2:0]
// FUNC -> I[5:3]
// ALUD -> I[8:6]
// RA -> A
// RB -> B
// H  -> mode32
// CI mux -> C0

// Status/Shifts:
// SHMUX -> I[9:6]
// STOPC -> I[5:0]
// CEM   -> ~nCEM
// CEN   -> ~nCEN
