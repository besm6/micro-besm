module testbench();

    // Input signals
    logic        clk;
    logic [63:0] word;
    logic        pe;
    logic        tkk;

    // Output signals
    logic  [3:0] ir;
    logic  [7:0] op;
    logic        extop;
    logic [19:0] addr;

    // Device under test
    decoder dut(word, pe, tkk,
        ir, op, extop, addr);

    // Status
    bit fail;

    // Read value from the variable.
    task verify(input check, input string message);
        if (!check) begin
            $display ("%s", message);
            fail = 1;
        end
    endtask

initial begin
$display("------------------------");
$dumpfile("test.vcd");
$dumpvars();
fail = 0;
clk = 0;

// ***************************************************
// * Test vectors for micro-BESM instruction decoder *
// ***************************************************
// 0000000000000000000000000000000000000000000000000000000000000001:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1
#2;

verify(ir === 'b0000, "Assert 0 : < ir !== 'b0000 >");	// Vector No: 0
verify(op === 'b00000000, "Assert 1 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000001:0:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 2
#2;

verify(ir === 'b0000, "Assert 4 : < ir !== 'b0000 >");	// Vector No: 1
verify(op === 'b00000000, "Assert 5 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 6 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 7 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000001:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 3
#2;

verify(ir === 'b0000, "Assert 8 : < ir !== 'b0000 >");	// Vector No: 2
verify(op === 'b00000000, "Assert 9 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 10 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 11 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000001:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 4
#2;

verify(ir === 'b0000, "Assert 12 : < ir !== 'b0000 >");	// Vector No: 3
verify(op === 'b00000000, "Assert 13 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 14 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 15 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000010:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 5
#2;

verify(ir === 'b0000, "Assert 16 : < ir !== 'b0000 >");	// Vector No: 4
verify(op === 'b00000000, "Assert 17 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 18 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 19 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000010:0:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 6
#2;

verify(ir === 'b0000, "Assert 20 : < ir !== 'b0000 >");	// Vector No: 5
verify(op === 'b00000000, "Assert 21 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 22 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 23 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000010:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 7
#2;

verify(ir === 'b0000, "Assert 24 : < ir !== 'b0000 >");	// Vector No: 6
verify(op === 'b00000000, "Assert 25 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 26 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 27 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000010:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 8
#2;

verify(ir === 'b0000, "Assert 28 : < ir !== 'b0000 >");	// Vector No: 7
verify(op === 'b00000000, "Assert 29 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 30 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 31 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000100:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 9
#2;

verify(ir === 'b0000, "Assert 32 : < ir !== 'b0000 >");	// Vector No: 8
verify(op === 'b00000000, "Assert 33 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 34 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 35 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000100:0:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 10
#2;

verify(ir === 'b0000, "Assert 36 : < ir !== 'b0000 >");	// Vector No: 9
verify(op === 'b00000000, "Assert 37 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 38 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 39 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000100:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 11
#2;

verify(ir === 'b0000, "Assert 40 : < ir !== 'b0000 >");	// Vector No: 10
verify(op === 'b00000000, "Assert 41 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 42 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 43 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000000100:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 12
#2;

verify(ir === 'b0000, "Assert 44 : < ir !== 'b0000 >");	// Vector No: 11
verify(op === 'b00000000, "Assert 45 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 46 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 47 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000001000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 13
#2;

verify(ir === 'b0000, "Assert 48 : < ir !== 'b0000 >");	// Vector No: 12
verify(op === 'b00000000, "Assert 49 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 50 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 51 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000001000:0:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 14
#2;

verify(ir === 'b0000, "Assert 52 : < ir !== 'b0000 >");	// Vector No: 13
verify(op === 'b00000000, "Assert 53 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 54 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 55 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000001000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 15
#2;

verify(ir === 'b0000, "Assert 56 : < ir !== 'b0000 >");	// Vector No: 14
verify(op === 'b00000000, "Assert 57 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 58 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 59 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000001000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 16
#2;

verify(ir === 'b0000, "Assert 60 : < ir !== 'b0000 >");	// Vector No: 15
verify(op === 'b00000000, "Assert 61 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 62 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 63 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000010000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 17
#2;

verify(ir === 'b0000, "Assert 64 : < ir !== 'b0000 >");	// Vector No: 16
verify(op === 'b00000000, "Assert 65 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 66 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 67 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000010000:0:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 18
#2;

verify(ir === 'b0000, "Assert 68 : < ir !== 'b0000 >");	// Vector No: 17
verify(op === 'b00000000, "Assert 69 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 70 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 71 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000010000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 19
#2;

verify(ir === 'b0000, "Assert 72 : < ir !== 'b0000 >");	// Vector No: 18
verify(op === 'b00000000, "Assert 73 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 74 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 75 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000010000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 20
#2;

verify(ir === 'b0000, "Assert 76 : < ir !== 'b0000 >");	// Vector No: 19
verify(op === 'b00000000, "Assert 77 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 78 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 79 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000100000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 21
#2;

verify(ir === 'b0000, "Assert 80 : < ir !== 'b0000 >");	// Vector No: 20
verify(op === 'b00000000, "Assert 81 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 82 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 83 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000100000:0:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 22
#2;

verify(ir === 'b0000, "Assert 84 : < ir !== 'b0000 >");	// Vector No: 21
verify(op === 'b00000000, "Assert 85 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 86 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 87 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000100000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 23
#2;

verify(ir === 'b0000, "Assert 88 : < ir !== 'b0000 >");	// Vector No: 22
verify(op === 'b00000000, "Assert 89 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 90 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 91 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000000100000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 24
#2;

verify(ir === 'b0000, "Assert 92 : < ir !== 'b0000 >");	// Vector No: 23
verify(op === 'b00000000, "Assert 93 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 94 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 95 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000001000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 25
#2;

verify(ir === 'b0000, "Assert 96 : < ir !== 'b0000 >");	// Vector No: 24
verify(op === 'b00000000, "Assert 97 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 98 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 99 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000001000000:0:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 26
#2;

verify(ir === 'b0000, "Assert 100 : < ir !== 'b0000 >");	// Vector No: 25
verify(op === 'b00000000, "Assert 101 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 102 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 103 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000001000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 27
#2;

verify(ir === 'b0000, "Assert 104 : < ir !== 'b0000 >");	// Vector No: 26
verify(op === 'b00000000, "Assert 105 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 106 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 107 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000001000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 28
#2;

verify(ir === 'b0000, "Assert 108 : < ir !== 'b0000 >");	// Vector No: 27
verify(op === 'b00000000, "Assert 109 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 110 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 111 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000010000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 29
#2;

verify(ir === 'b0000, "Assert 112 : < ir !== 'b0000 >");	// Vector No: 28
verify(op === 'b00000000, "Assert 113 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 114 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 115 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000010000000:0:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 30
#2;

verify(ir === 'b0000, "Assert 116 : < ir !== 'b0000 >");	// Vector No: 29
verify(op === 'b00000000, "Assert 117 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 118 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 119 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000010000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 31
#2;

verify(ir === 'b0000, "Assert 120 : < ir !== 'b0000 >");	// Vector No: 30
verify(op === 'b00000000, "Assert 121 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 122 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 123 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000010000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 32
#2;

verify(ir === 'b0000, "Assert 124 : < ir !== 'b0000 >");	// Vector No: 31
verify(op === 'b00000000, "Assert 125 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 126 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 127 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000100000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 33
#2;

verify(ir === 'b0000, "Assert 128 : < ir !== 'b0000 >");	// Vector No: 32
verify(op === 'b00000000, "Assert 129 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 130 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 131 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000100000000:0:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 34
#2;

verify(ir === 'b0000, "Assert 132 : < ir !== 'b0000 >");	// Vector No: 33
verify(op === 'b00000000, "Assert 133 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 134 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 135 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000100000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 35
#2;

verify(ir === 'b0000, "Assert 136 : < ir !== 'b0000 >");	// Vector No: 34
verify(op === 'b00000000, "Assert 137 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 138 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 139 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000000100000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 36
#2;

verify(ir === 'b0000, "Assert 140 : < ir !== 'b0000 >");	// Vector No: 35
verify(op === 'b00000000, "Assert 141 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 142 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 143 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000001000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 37
#2;

verify(ir === 'b0000, "Assert 144 : < ir !== 'b0000 >");	// Vector No: 36
verify(op === 'b00000000, "Assert 145 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 146 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 147 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000001000000000:0:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 38
#2;

verify(ir === 'b0000, "Assert 148 : < ir !== 'b0000 >");	// Vector No: 37
verify(op === 'b00000000, "Assert 149 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 150 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 151 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000001000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 39
#2;

verify(ir === 'b0000, "Assert 152 : < ir !== 'b0000 >");	// Vector No: 38
verify(op === 'b00000000, "Assert 153 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 154 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 155 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000001000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 40
#2;

verify(ir === 'b0000, "Assert 156 : < ir !== 'b0000 >");	// Vector No: 39
verify(op === 'b00000000, "Assert 157 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 158 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 159 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000010000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 41
#2;

verify(ir === 'b0000, "Assert 160 : < ir !== 'b0000 >");	// Vector No: 40
verify(op === 'b00000000, "Assert 161 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 162 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 163 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000010000000000:0:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 42
#2;

verify(ir === 'b0000, "Assert 164 : < ir !== 'b0000 >");	// Vector No: 41
verify(op === 'b00000000, "Assert 165 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 166 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 167 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000010000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 43
#2;

verify(ir === 'b0000, "Assert 168 : < ir !== 'b0000 >");	// Vector No: 42
verify(op === 'b00000000, "Assert 169 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 170 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 171 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000010000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 44
#2;

verify(ir === 'b0000, "Assert 172 : < ir !== 'b0000 >");	// Vector No: 43
verify(op === 'b00000000, "Assert 173 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 174 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 175 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000100000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 45
#2;

verify(ir === 'b0000, "Assert 176 : < ir !== 'b0000 >");	// Vector No: 44
verify(op === 'b00000000, "Assert 177 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 178 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 179 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000100000000000:0:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 46
#2;

verify(ir === 'b0000, "Assert 180 : < ir !== 'b0000 >");	// Vector No: 45
verify(op === 'b00000000, "Assert 181 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 182 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 183 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000100000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 47
#2;

verify(ir === 'b0000, "Assert 184 : < ir !== 'b0000 >");	// Vector No: 46
verify(op === 'b00000000, "Assert 185 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 186 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 187 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000000100000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 48
#2;

verify(ir === 'b0000, "Assert 188 : < ir !== 'b0000 >");	// Vector No: 47
verify(op === 'b00000000, "Assert 189 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 190 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 191 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000001000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 49
#2;

verify(ir === 'b0000, "Assert 192 : < ir !== 'b0000 >");	// Vector No: 48
verify(op === 'b00000000, "Assert 193 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 194 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 195 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000001000000000000:0:1:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 50
#2;

verify(ir === 'b0000, "Assert 196 : < ir !== 'b0000 >");	// Vector No: 49
verify(op === 'b00000000, "Assert 197 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 198 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 199 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000001000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 51
#2;

verify(ir === 'b0000, "Assert 200 : < ir !== 'b0000 >");	// Vector No: 50
verify(op === 'b00000000, "Assert 201 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 202 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 203 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000001000000000000:1:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 52
#2;

verify(ir === 'b0000, "Assert 204 : < ir !== 'b0000 >");	// Vector No: 51
verify(op === 'b00000000, "Assert 205 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 206 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 207 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000010000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 53
#2;

verify(ir === 'b0000, "Assert 208 : < ir !== 'b0000 >");	// Vector No: 52
verify(op === 'b00000000, "Assert 209 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 210 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 211 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000010000000000000:0:1:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 54
#2;

verify(ir === 'b0000, "Assert 212 : < ir !== 'b0000 >");	// Vector No: 53
verify(op === 'b00000000, "Assert 213 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 214 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 215 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000010000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 55
#2;

verify(ir === 'b0000, "Assert 216 : < ir !== 'b0000 >");	// Vector No: 54
verify(op === 'b00000000, "Assert 217 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 218 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 219 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000010000000000000:1:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 56
#2;

verify(ir === 'b0000, "Assert 220 : < ir !== 'b0000 >");	// Vector No: 55
verify(op === 'b00000000, "Assert 221 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 222 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 223 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000100000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 57
#2;

verify(ir === 'b0000, "Assert 224 : < ir !== 'b0000 >");	// Vector No: 56
verify(op === 'b00000000, "Assert 225 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 226 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 227 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000100000000000000:0:1:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 58
#2;

verify(ir === 'b0000, "Assert 228 : < ir !== 'b0000 >");	// Vector No: 57
verify(op === 'b00000000, "Assert 229 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 230 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 231 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000100000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 59
#2;

verify(ir === 'b0000, "Assert 232 : < ir !== 'b0000 >");	// Vector No: 58
verify(op === 'b00000000, "Assert 233 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 234 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 235 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000000100000000000000:1:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 60
#2;

verify(ir === 'b0000, "Assert 236 : < ir !== 'b0000 >");	// Vector No: 59
verify(op === 'b00000000, "Assert 237 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 238 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 239 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000001000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 61
#2;

verify(ir === 'b0000, "Assert 240 : < ir !== 'b0000 >");	// Vector No: 60
verify(op === 'b00000000, "Assert 241 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 242 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 243 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000001000000000000000:0:1:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 62
#2;

verify(ir === 'b0000, "Assert 244 : < ir !== 'b0000 >");	// Vector No: 61
verify(op === 'b00000000, "Assert 245 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 246 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 247 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000001000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 63
#2;

verify(ir === 'b0000, "Assert 248 : < ir !== 'b0000 >");	// Vector No: 62
verify(op === 'b00000000, "Assert 249 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 250 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 251 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000001000000000000000:1:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 64
#2;

verify(ir === 'b0000, "Assert 252 : < ir !== 'b0000 >");	// Vector No: 63
verify(op === 'b00000000, "Assert 253 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 254 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 255 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000010000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 65
#2;

verify(ir === 'b0000, "Assert 256 : < ir !== 'b0000 >");	// Vector No: 64
verify(op === 'b00000000, "Assert 257 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 258 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 259 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000010000000000000000:0:1:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 66
#2;

verify(ir === 'b0000, "Assert 260 : < ir !== 'b0000 >");	// Vector No: 65
verify(op === 'b00000000, "Assert 261 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 262 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 263 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000010000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 67
#2;

verify(ir === 'b0000, "Assert 264 : < ir !== 'b0000 >");	// Vector No: 66
verify(op === 'b00000000, "Assert 265 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 266 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 267 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000010000000000000000:1:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 68
#2;

verify(ir === 'b0000, "Assert 268 : < ir !== 'b0000 >");	// Vector No: 67
verify(op === 'b00000000, "Assert 269 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 270 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 271 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000100000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 69
#2;

verify(ir === 'b0000, "Assert 272 : < ir !== 'b0000 >");	// Vector No: 68
verify(op === 'b00000000, "Assert 273 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 274 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 275 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000100000000000000000:0:1:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 70
#2;

verify(ir === 'b0000, "Assert 276 : < ir !== 'b0000 >");	// Vector No: 69
verify(op === 'b00000000, "Assert 277 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 278 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 279 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000100000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 71
#2;

verify(ir === 'b0000, "Assert 280 : < ir !== 'b0000 >");	// Vector No: 70
verify(op === 'b00000000, "Assert 281 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 282 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 283 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000000100000000000000000:1:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 72
#2;

verify(ir === 'b0000, "Assert 284 : < ir !== 'b0000 >");	// Vector No: 71
verify(op === 'b00000000, "Assert 285 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 286 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 287 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000001000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 73
#2;

verify(ir === 'b0000, "Assert 288 : < ir !== 'b0000 >");	// Vector No: 72
verify(op === 'b00000000, "Assert 289 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 290 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 291 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000001000000000000000000:0:1:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 74
#2;

verify(ir === 'b0000, "Assert 292 : < ir !== 'b0000 >");	// Vector No: 73
verify(op === 'b00000000, "Assert 293 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 294 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 295 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000001000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 75
#2;

verify(ir === 'b0000, "Assert 296 : < ir !== 'b0000 >");	// Vector No: 74
verify(op === 'b00000000, "Assert 297 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 298 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 299 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000001000000000000000000:1:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 76
#2;

verify(ir === 'b0000, "Assert 300 : < ir !== 'b0000 >");	// Vector No: 75
verify(op === 'b00000000, "Assert 301 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 302 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 303 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000010000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 77
#2;

verify(ir === 'b0000, "Assert 304 : < ir !== 'b0000 >");	// Vector No: 76
verify(op === 'b00000000, "Assert 305 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 306 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 307 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000010000000000000000000:0:1:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 78
#2;

verify(ir === 'b0000, "Assert 308 : < ir !== 'b0000 >");	// Vector No: 77
verify(op === 'b00000000, "Assert 309 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 310 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 311 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000010000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 79
#2;

verify(ir === 'b0000, "Assert 312 : < ir !== 'b0000 >");	// Vector No: 78
verify(op === 'b00000000, "Assert 313 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 314 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 315 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000010000000000000000000:1:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 80
#2;

verify(ir === 'b0000, "Assert 316 : < ir !== 'b0000 >");	// Vector No: 79
verify(op === 'b00000000, "Assert 317 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 318 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 319 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 81
#2;

verify(ir === 'b0000, "Assert 320 : < ir !== 'b0000 >");	// Vector No: 80
verify(op === 'b00000000, "Assert 321 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 322 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 323 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000100000000000000000000:0:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 82
#2;

verify(ir === 'b0000, "Assert 324 : < ir !== 'b0000 >");	// Vector No: 81
verify(op === 'b00000001, "Assert 325 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 326 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 327 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 83
#2;

verify(ir === 'b0000, "Assert 328 : < ir !== 'b0000 >");	// Vector No: 82
verify(op === 'b00000000, "Assert 329 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 330 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 331 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000000100000000000000000000:1:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 84
#2;

verify(ir === 'b0000, "Assert 332 : < ir !== 'b0000 >");	// Vector No: 83
verify(op === 'b00000000, "Assert 333 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 334 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 335 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000001000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 85
#2;

verify(ir === 'b0000, "Assert 336 : < ir !== 'b0000 >");	// Vector No: 84
verify(op === 'b00000000, "Assert 337 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 338 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 339 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000001000000000000000000000:0:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 86
#2;

verify(ir === 'b0000, "Assert 340 : < ir !== 'b0000 >");	// Vector No: 85
verify(op === 'b00000010, "Assert 341 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 342 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 343 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000001000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 87
#2;

verify(ir === 'b0000, "Assert 344 : < ir !== 'b0000 >");	// Vector No: 86
verify(op === 'b00000000, "Assert 345 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 346 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 347 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000001000000000000000000000:1:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 88
#2;

verify(ir === 'b0000, "Assert 348 : < ir !== 'b0000 >");	// Vector No: 87
verify(op === 'b00000000, "Assert 349 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 350 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 351 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000010000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 89
#2;

verify(ir === 'b0000, "Assert 352 : < ir !== 'b0000 >");	// Vector No: 88
verify(op === 'b00000000, "Assert 353 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 354 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 355 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000010000000000000000000000:0:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 90
#2;

verify(ir === 'b0000, "Assert 356 : < ir !== 'b0000 >");	// Vector No: 89
verify(op === 'b00000100, "Assert 357 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 358 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 359 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000010000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 91
#2;

verify(ir === 'b0000, "Assert 360 : < ir !== 'b0000 >");	// Vector No: 90
verify(op === 'b00000000, "Assert 361 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 362 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 363 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000010000000000000000000000:1:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 92
#2;

verify(ir === 'b0000, "Assert 364 : < ir !== 'b0000 >");	// Vector No: 91
verify(op === 'b00000000, "Assert 365 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 366 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 367 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000100000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 93
#2;

verify(ir === 'b0000, "Assert 368 : < ir !== 'b0000 >");	// Vector No: 92
verify(op === 'b00000000, "Assert 369 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 370 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 371 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000100000000000000000000000:0:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 94
#2;

verify(ir === 'b0000, "Assert 372 : < ir !== 'b0000 >");	// Vector No: 93
verify(op === 'b00001000, "Assert 373 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 374 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 375 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000100000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 95
#2;

verify(ir === 'b0000, "Assert 376 : < ir !== 'b0000 >");	// Vector No: 94
verify(op === 'b00000000, "Assert 377 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 378 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 379 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000000100000000000000000000000:1:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 96
#2;

verify(ir === 'b0000, "Assert 380 : < ir !== 'b0000 >");	// Vector No: 95
verify(op === 'b00000000, "Assert 381 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 382 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 383 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000001000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 97
#2;

verify(ir === 'b0000, "Assert 384 : < ir !== 'b0000 >");	// Vector No: 96
verify(op === 'b00000000, "Assert 385 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 386 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 387 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000001000000000000000000000000:0:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 98
#2;

verify(ir === 'b0000, "Assert 388 : < ir !== 'b0000 >");	// Vector No: 97
verify(op === 'b00010000, "Assert 389 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 390 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 391 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000001000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 99
#2;

verify(ir === 'b0000, "Assert 392 : < ir !== 'b0000 >");	// Vector No: 98
verify(op === 'b00000000, "Assert 393 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 394 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 395 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000001000000000000000000000000:1:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 100
#2;

verify(ir === 'b0000, "Assert 396 : < ir !== 'b0000 >");	// Vector No: 99
verify(op === 'b00000001, "Assert 397 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 398 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 399 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000010000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 101
#2;

verify(ir === 'b0000, "Assert 400 : < ir !== 'b0000 >");	// Vector No: 100
verify(op === 'b00000000, "Assert 401 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 402 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 403 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000010000000000000000000000000:0:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 102
#2;

verify(ir === 'b0000, "Assert 404 : < ir !== 'b0000 >");	// Vector No: 101
verify(op === 'b00100000, "Assert 405 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 406 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 407 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000010000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 103
#2;

verify(ir === 'b0000, "Assert 408 : < ir !== 'b0000 >");	// Vector No: 102
verify(op === 'b00000000, "Assert 409 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 410 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 411 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000010000000000000000000000000:1:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 104
#2;

verify(ir === 'b0000, "Assert 412 : < ir !== 'b0000 >");	// Vector No: 103
verify(op === 'b00000010, "Assert 413 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 414 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 415 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000100000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 105
#2;

verify(ir === 'b0000, "Assert 416 : < ir !== 'b0000 >");	// Vector No: 104
verify(op === 'b00000000, "Assert 417 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 418 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 419 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000100000000000000000000000000:0:1:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 106
#2;

verify(ir === 'b0000, "Assert 420 : < ir !== 'b0000 >");	// Vector No: 105
verify(op === 'b01000000, "Assert 421 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 422 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 423 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000100000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 107
#2;

verify(ir === 'b0000, "Assert 424 : < ir !== 'b0000 >");	// Vector No: 106
verify(op === 'b00000000, "Assert 425 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 426 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 427 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000100000000000000000000000000:1:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 108
#2;

verify(ir === 'b0000, "Assert 428 : < ir !== 'b0000 >");	// Vector No: 107
verify(op === 'b00000100, "Assert 429 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 430 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 431 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000001000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 109
#2;

verify(ir === 'b0000, "Assert 432 : < ir !== 'b0000 >");	// Vector No: 108
verify(op === 'b00000000, "Assert 433 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 434 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 435 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000001000000000000000000000000000:0:1:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 110
#2;

verify(ir === 'b0000, "Assert 436 : < ir !== 'b0000 >");	// Vector No: 109
verify(op === 'b10000000, "Assert 437 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 438 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 439 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000001000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 111
#2;

verify(ir === 'b0000, "Assert 440 : < ir !== 'b0000 >");	// Vector No: 110
verify(op === 'b00000000, "Assert 441 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 442 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 443 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000001000000000000000000000000000:1:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 112
#2;

verify(ir === 'b0000, "Assert 444 : < ir !== 'b0000 >");	// Vector No: 111
verify(op === 'b00001000, "Assert 445 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 446 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 447 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 113
#2;

verify(ir === 'b0000, "Assert 448 : < ir !== 'b0000 >");	// Vector No: 112
verify(op === 'b00000000, "Assert 449 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 450 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 451 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010000000000000000000000000000:0:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 114
#2;

verify(ir === 'b0001, "Assert 452 : < ir !== 'b0001 >");	// Vector No: 113
verify(op === 'b00000000, "Assert 453 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 454 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 455 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 115
#2;

verify(ir === 'b0000, "Assert 456 : < ir !== 'b0000 >");	// Vector No: 114
verify(op === 'b00000000, "Assert 457 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 458 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 459 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010000000000000000000000000000:1:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 116
#2;

verify(ir === 'b0000, "Assert 460 : < ir !== 'b0000 >");	// Vector No: 115
verify(op === 'b00010000, "Assert 461 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 462 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 463 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 117
#2;

verify(ir === 'b0000, "Assert 464 : < ir !== 'b0000 >");	// Vector No: 116
verify(op === 'b00000000, "Assert 465 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 466 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 467 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100000000000000000000000000000:0:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 118
#2;

verify(ir === 'b0010, "Assert 468 : < ir !== 'b0010 >");	// Vector No: 117
verify(op === 'b00000000, "Assert 469 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 470 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 471 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 119
#2;

verify(ir === 'b0000, "Assert 472 : < ir !== 'b0000 >");	// Vector No: 118
verify(op === 'b00000000, "Assert 473 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 474 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 475 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100000000000000000000000000000:1:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 120
#2;

verify(ir === 'b0000, "Assert 476 : < ir !== 'b0000 >");	// Vector No: 119
verify(op === 'b00100000, "Assert 477 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 478 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 479 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 121
#2;

verify(ir === 'b0000, "Assert 480 : < ir !== 'b0000 >");	// Vector No: 120
verify(op === 'b00000000, "Assert 481 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 482 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 483 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000000000000000000000000000000:0:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 122
#2;

verify(ir === 'b0100, "Assert 484 : < ir !== 'b0100 >");	// Vector No: 121
verify(op === 'b00000000, "Assert 485 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 486 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 487 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 123
#2;

verify(ir === 'b0000, "Assert 488 : < ir !== 'b0000 >");	// Vector No: 122
verify(op === 'b00000000, "Assert 489 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 490 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 491 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000000000000000000000000000000:1:1:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 124
#2;

verify(ir === 'b0000, "Assert 492 : < ir !== 'b0000 >");	// Vector No: 123
verify(op === 'b01000000, "Assert 493 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 494 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 495 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 125
#2;

verify(ir === 'b0000, "Assert 496 : < ir !== 'b0000 >");	// Vector No: 124
verify(op === 'b00000000, "Assert 497 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 498 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 499 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 126
#2;

verify(ir === 'b1000, "Assert 500 : < ir !== 'b1000 >");	// Vector No: 125
verify(op === 'b00000000, "Assert 501 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 502 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 503 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 127
#2;

verify(ir === 'b0000, "Assert 504 : < ir !== 'b0000 >");	// Vector No: 126
verify(op === 'b00000000, "Assert 505 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 506 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 507 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 128
#2;

verify(ir === 'b0000, "Assert 508 : < ir !== 'b0000 >");	// Vector No: 127
verify(op === 'b00000000, "Assert 509 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 510 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 511 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 129
#2;

verify(ir === 'b0000, "Assert 512 : < ir !== 'b0000 >");	// Vector No: 128
verify(op === 'b00000000, "Assert 513 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 514 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 515 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 130
#2;

verify(ir === 'b0000, "Assert 516 : < ir !== 'b0000 >");	// Vector No: 129
verify(op === 'b00000000, "Assert 517 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 518 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 519 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 131
#2;

verify(ir === 'b0000, "Assert 520 : < ir !== 'b0000 >");	// Vector No: 130
verify(op === 'b00000000, "Assert 521 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 522 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 523 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000000000000000000000000000000:1:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 132
#2;

verify(ir === 'b0001, "Assert 524 : < ir !== 'b0001 >");	// Vector No: 131
verify(op === 'b00000000, "Assert 525 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 526 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 527 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 133
#2;

verify(ir === 'b0000, "Assert 528 : < ir !== 'b0000 >");	// Vector No: 132
verify(op === 'b00000000, "Assert 529 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 530 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 531 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 134
#2;

verify(ir === 'b0000, "Assert 532 : < ir !== 'b0000 >");	// Vector No: 133
verify(op === 'b00000000, "Assert 533 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 534 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 535 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 135
#2;

verify(ir === 'b0000, "Assert 536 : < ir !== 'b0000 >");	// Vector No: 134
verify(op === 'b00000000, "Assert 537 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 538 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 539 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000000000000000000000000000000:1:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 136
#2;

verify(ir === 'b0010, "Assert 540 : < ir !== 'b0010 >");	// Vector No: 135
verify(op === 'b00000000, "Assert 541 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 542 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 543 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 137
#2;

verify(ir === 'b0000, "Assert 544 : < ir !== 'b0000 >");	// Vector No: 136
verify(op === 'b00000000, "Assert 545 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 546 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 547 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 138
#2;

verify(ir === 'b0000, "Assert 548 : < ir !== 'b0000 >");	// Vector No: 137
verify(op === 'b00000000, "Assert 549 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 550 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 551 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 139
#2;

verify(ir === 'b0000, "Assert 552 : < ir !== 'b0000 >");	// Vector No: 138
verify(op === 'b00000000, "Assert 553 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 554 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 555 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000000000000000000000000000000:1:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 140
#2;

verify(ir === 'b0100, "Assert 556 : < ir !== 'b0100 >");	// Vector No: 139
verify(op === 'b00000000, "Assert 557 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 558 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 559 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000000000000000000000000000000:0:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 141
#2;

verify(ir === 'b0000, "Assert 560 : < ir !== 'b0000 >");	// Vector No: 140
verify(op === 'b00000000, "Assert 561 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 562 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 563 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 142
#2;

verify(ir === 'b0000, "Assert 564 : < ir !== 'b0000 >");	// Vector No: 141
verify(op === 'b00000000, "Assert 565 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 566 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 567 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 143
#2;

verify(ir === 'b0000, "Assert 568 : < ir !== 'b0000 >");	// Vector No: 142
verify(op === 'b00000000, "Assert 569 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 570 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 571 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000000000000000000000000000000:1:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 144
#2;

verify(ir === 'b1000, "Assert 572 : < ir !== 'b1000 >");	// Vector No: 143
verify(op === 'b00000000, "Assert 573 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 574 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 575 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000000000000000000000000000000:0:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 145
#2;

verify(ir === 'b0000, "Assert 576 : < ir !== 'b0000 >");	// Vector No: 144
verify(op === 'b00000000, "Assert 577 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 578 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 579 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 146
#2;

verify(ir === 'b0000, "Assert 580 : < ir !== 'b0000 >");	// Vector No: 145
verify(op === 'b00000000, "Assert 581 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 582 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 583 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 147
#2;

verify(ir === 'b0000, "Assert 584 : < ir !== 'b0000 >");	// Vector No: 146
verify(op === 'b00000000, "Assert 585 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 586 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 587 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 148
#2;

verify(ir === 'b0000, "Assert 588 : < ir !== 'b0000 >");	// Vector No: 147
verify(op === 'b00000000, "Assert 589 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 590 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 591 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000000000000000000000000000000:0:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 149
#2;

verify(ir === 'b0000, "Assert 592 : < ir !== 'b0000 >");	// Vector No: 148
verify(op === 'b00000000, "Assert 593 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 594 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 595 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 150
#2;

verify(ir === 'b0000, "Assert 596 : < ir !== 'b0000 >");	// Vector No: 149
verify(op === 'b00000000, "Assert 597 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 598 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 599 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 151
#2;

verify(ir === 'b0000, "Assert 600 : < ir !== 'b0000 >");	// Vector No: 150
verify(op === 'b00000000, "Assert 601 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 602 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 603 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 152
#2;

verify(ir === 'b0000, "Assert 604 : < ir !== 'b0000 >");	// Vector No: 151
verify(op === 'b00000000, "Assert 605 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 606 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 607 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000000000000000000000000000000:0:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 153
#2;

verify(ir === 'b0000, "Assert 608 : < ir !== 'b0000 >");	// Vector No: 152
verify(op === 'b00000000, "Assert 609 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 610 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 611 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 154
#2;

verify(ir === 'b0000, "Assert 612 : < ir !== 'b0000 >");	// Vector No: 153
verify(op === 'b00000000, "Assert 613 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 614 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 615 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 155
#2;

verify(ir === 'b0000, "Assert 616 : < ir !== 'b0000 >");	// Vector No: 154
verify(op === 'b00000000, "Assert 617 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 618 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 619 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 156
#2;

verify(ir === 'b0000, "Assert 620 : < ir !== 'b0000 >");	// Vector No: 155
verify(op === 'b00000000, "Assert 621 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 622 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 623 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000000000000000000000000000000:0:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 157
#2;

verify(ir === 'b0000, "Assert 624 : < ir !== 'b0000 >");	// Vector No: 156
verify(op === 'b00000000, "Assert 625 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 626 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 627 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 158
#2;

verify(ir === 'b0000, "Assert 628 : < ir !== 'b0000 >");	// Vector No: 157
verify(op === 'b00000000, "Assert 629 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 630 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 631 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 159
#2;

verify(ir === 'b0000, "Assert 632 : < ir !== 'b0000 >");	// Vector No: 158
verify(op === 'b00000000, "Assert 633 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 634 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 635 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 160
#2;

verify(ir === 'b0000, "Assert 636 : < ir !== 'b0000 >");	// Vector No: 159
verify(op === 'b00000000, "Assert 637 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 638 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 639 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000000000000000000000000000000:0:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 161
#2;

verify(ir === 'b0000, "Assert 640 : < ir !== 'b0000 >");	// Vector No: 160
verify(op === 'b00000000, "Assert 641 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 642 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 643 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 162
#2;

verify(ir === 'b0000, "Assert 644 : < ir !== 'b0000 >");	// Vector No: 161
verify(op === 'b00000000, "Assert 645 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 646 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 647 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 163
#2;

verify(ir === 'b0000, "Assert 648 : < ir !== 'b0000 >");	// Vector No: 162
verify(op === 'b00000000, "Assert 649 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 650 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 651 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 164
#2;

verify(ir === 'b0000, "Assert 652 : < ir !== 'b0000 >");	// Vector No: 163
verify(op === 'b00000000, "Assert 653 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 654 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 655 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000000000000000000000000000000:0:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 165
#2;

verify(ir === 'b0000, "Assert 656 : < ir !== 'b0000 >");	// Vector No: 164
verify(op === 'b00000000, "Assert 657 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 658 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 659 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 166
#2;

verify(ir === 'b0000, "Assert 660 : < ir !== 'b0000 >");	// Vector No: 165
verify(op === 'b00000000, "Assert 661 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 662 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 663 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 167
#2;

verify(ir === 'b0000, "Assert 664 : < ir !== 'b0000 >");	// Vector No: 166
verify(op === 'b00000000, "Assert 665 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 666 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 667 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 168
#2;

verify(ir === 'b0000, "Assert 668 : < ir !== 'b0000 >");	// Vector No: 167
verify(op === 'b00000000, "Assert 669 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 670 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 671 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000000000000000000000000000000:0:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 169
#2;

verify(ir === 'b0000, "Assert 672 : < ir !== 'b0000 >");	// Vector No: 168
verify(op === 'b00000000, "Assert 673 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 674 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 675 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 170
#2;

verify(ir === 'b0000, "Assert 676 : < ir !== 'b0000 >");	// Vector No: 169
verify(op === 'b00000000, "Assert 677 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 678 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 679 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 171
#2;

verify(ir === 'b0000, "Assert 680 : < ir !== 'b0000 >");	// Vector No: 170
verify(op === 'b00000000, "Assert 681 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 682 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 683 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 172
#2;

verify(ir === 'b0000, "Assert 684 : < ir !== 'b0000 >");	// Vector No: 171
verify(op === 'b00000000, "Assert 685 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 686 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 687 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000000000000000000000000000000:0:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 173
#2;

verify(ir === 'b0000, "Assert 688 : < ir !== 'b0000 >");	// Vector No: 172
verify(op === 'b00000000, "Assert 689 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 690 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 691 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 174
#2;

verify(ir === 'b0000, "Assert 692 : < ir !== 'b0000 >");	// Vector No: 173
verify(op === 'b00000000, "Assert 693 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 694 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 695 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 175
#2;

verify(ir === 'b0000, "Assert 696 : < ir !== 'b0000 >");	// Vector No: 174
verify(op === 'b00000000, "Assert 697 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 698 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 699 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 176
#2;

verify(ir === 'b0000, "Assert 700 : < ir !== 'b0000 >");	// Vector No: 175
verify(op === 'b00000000, "Assert 701 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 702 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 703 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000000000000000000000000000000:0:0:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 177
#2;

verify(ir === 'b0000, "Assert 704 : < ir !== 'b0000 >");	// Vector No: 176
verify(op === 'b00000000, "Assert 705 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 706 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 707 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 178
#2;

verify(ir === 'b0000, "Assert 708 : < ir !== 'b0000 >");	// Vector No: 177
verify(op === 'b00000000, "Assert 709 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 710 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 711 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 179
#2;

verify(ir === 'b0000, "Assert 712 : < ir !== 'b0000 >");	// Vector No: 178
verify(op === 'b00000000, "Assert 713 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 714 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 715 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 180
#2;

verify(ir === 'b0000, "Assert 716 : < ir !== 'b0000 >");	// Vector No: 179
verify(op === 'b00000000, "Assert 717 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 718 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 719 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000000000000000000000000000000:0:0:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 181
#2;

verify(ir === 'b0000, "Assert 720 : < ir !== 'b0000 >");	// Vector No: 180
verify(op === 'b00000000, "Assert 721 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 722 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 723 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 182
#2;

verify(ir === 'b0000, "Assert 724 : < ir !== 'b0000 >");	// Vector No: 181
verify(op === 'b00000000, "Assert 725 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 726 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 727 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 183
#2;

verify(ir === 'b0000, "Assert 728 : < ir !== 'b0000 >");	// Vector No: 182
verify(op === 'b00000000, "Assert 729 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 730 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 731 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 184
#2;

verify(ir === 'b0000, "Assert 732 : < ir !== 'b0000 >");	// Vector No: 183
verify(op === 'b00000000, "Assert 733 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 734 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 735 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000000000000000000000000000000:0:0:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 185
#2;

verify(ir === 'b0000, "Assert 736 : < ir !== 'b0000 >");	// Vector No: 184
verify(op === 'b00000000, "Assert 737 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 738 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 739 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 186
#2;

verify(ir === 'b0000, "Assert 740 : < ir !== 'b0000 >");	// Vector No: 185
verify(op === 'b00000000, "Assert 741 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 742 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 743 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 187
#2;

verify(ir === 'b0000, "Assert 744 : < ir !== 'b0000 >");	// Vector No: 186
verify(op === 'b00000000, "Assert 745 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 746 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 747 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 188
#2;

verify(ir === 'b0000, "Assert 748 : < ir !== 'b0000 >");	// Vector No: 187
verify(op === 'b00000000, "Assert 749 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 750 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 751 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000000000000000000000000000000:0:0:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 189
#2;

verify(ir === 'b0000, "Assert 752 : < ir !== 'b0000 >");	// Vector No: 188
verify(op === 'b00000000, "Assert 753 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 754 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 755 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 190
#2;

verify(ir === 'b0000, "Assert 756 : < ir !== 'b0000 >");	// Vector No: 189
verify(op === 'b00000000, "Assert 757 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 758 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 759 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 191
#2;

verify(ir === 'b0000, "Assert 760 : < ir !== 'b0000 >");	// Vector No: 190
verify(op === 'b00000000, "Assert 761 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 762 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 763 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 192
#2;

verify(ir === 'b0000, "Assert 764 : < ir !== 'b0000 >");	// Vector No: 191
verify(op === 'b00000000, "Assert 765 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 766 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 767 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000000000000000000000000000000:0:0:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 193
#2;

verify(ir === 'b0000, "Assert 768 : < ir !== 'b0000 >");	// Vector No: 192
verify(op === 'b00000000, "Assert 769 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 770 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 771 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 194
#2;

verify(ir === 'b0000, "Assert 772 : < ir !== 'b0000 >");	// Vector No: 193
verify(op === 'b00000000, "Assert 773 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 774 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 775 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000000000000000000000000000000:1:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 195
#2;

verify(ir === 'b0000, "Assert 776 : < ir !== 'b0000 >");	// Vector No: 194
verify(op === 'b00000001, "Assert 777 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 778 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 779 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 196
#2;

verify(ir === 'b0000, "Assert 780 : < ir !== 'b0000 >");	// Vector No: 195
verify(op === 'b00000000, "Assert 781 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 782 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 783 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000000000000000000000000000000:0:0:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 197
#2;

verify(ir === 'b0000, "Assert 784 : < ir !== 'b0000 >");	// Vector No: 196
verify(op === 'b00000000, "Assert 785 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 786 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 787 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 198
#2;

verify(ir === 'b0000, "Assert 788 : < ir !== 'b0000 >");	// Vector No: 197
verify(op === 'b00000000, "Assert 789 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 790 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 791 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000000000000000000000000000000:1:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 199
#2;

verify(ir === 'b0000, "Assert 792 : < ir !== 'b0000 >");	// Vector No: 198
verify(op === 'b00000010, "Assert 793 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 794 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 795 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 200
#2;

verify(ir === 'b0000, "Assert 796 : < ir !== 'b0000 >");	// Vector No: 199
verify(op === 'b00000000, "Assert 797 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 798 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 799 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000000000000000000000000000000:0:0:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 201
#2;

verify(ir === 'b0000, "Assert 800 : < ir !== 'b0000 >");	// Vector No: 200
verify(op === 'b00000000, "Assert 801 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 802 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 803 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 202
#2;

verify(ir === 'b0000, "Assert 804 : < ir !== 'b0000 >");	// Vector No: 201
verify(op === 'b00000000, "Assert 805 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 806 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 807 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000000000000000000000000000000:1:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 203
#2;

verify(ir === 'b0000, "Assert 808 : < ir !== 'b0000 >");	// Vector No: 202
verify(op === 'b00000100, "Assert 809 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 810 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 811 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 204
#2;

verify(ir === 'b0000, "Assert 812 : < ir !== 'b0000 >");	// Vector No: 203
verify(op === 'b00000000, "Assert 813 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 814 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 815 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000000000000000000000000000000:0:0:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 205
#2;

verify(ir === 'b0000, "Assert 816 : < ir !== 'b0000 >");	// Vector No: 204
verify(op === 'b00000000, "Assert 817 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 818 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 819 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 206
#2;

verify(ir === 'b0000, "Assert 820 : < ir !== 'b0000 >");	// Vector No: 205
verify(op === 'b00000000, "Assert 821 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 822 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 823 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000000000000000000000000000000:1:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 207
#2;

verify(ir === 'b0000, "Assert 824 : < ir !== 'b0000 >");	// Vector No: 206
verify(op === 'b00001000, "Assert 825 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 826 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 827 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 208
#2;

verify(ir === 'b0000, "Assert 828 : < ir !== 'b0000 >");	// Vector No: 207
verify(op === 'b00000000, "Assert 829 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 830 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 831 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000000000000000000000000000000:0:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 209
#2;

verify(ir === 'b0000, "Assert 832 : < ir !== 'b0000 >");	// Vector No: 208
verify(op === 'b00000001, "Assert 833 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 834 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 835 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 210
#2;

verify(ir === 'b0000, "Assert 836 : < ir !== 'b0000 >");	// Vector No: 209
verify(op === 'b00000000, "Assert 837 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 838 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 839 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000000000000000000000000000000:1:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 211
#2;

verify(ir === 'b0000, "Assert 840 : < ir !== 'b0000 >");	// Vector No: 210
verify(op === 'b00010000, "Assert 841 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 842 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 843 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 212
#2;

verify(ir === 'b0000, "Assert 844 : < ir !== 'b0000 >");	// Vector No: 211
verify(op === 'b00000000, "Assert 845 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 846 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 847 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000000000000000000000000000000:0:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 213
#2;

verify(ir === 'b0000, "Assert 848 : < ir !== 'b0000 >");	// Vector No: 212
verify(op === 'b00000010, "Assert 849 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 850 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 851 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 214
#2;

verify(ir === 'b0000, "Assert 852 : < ir !== 'b0000 >");	// Vector No: 213
verify(op === 'b00000000, "Assert 853 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 854 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 855 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000000000000000000000000000000:1:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 215
#2;

verify(ir === 'b0000, "Assert 856 : < ir !== 'b0000 >");	// Vector No: 214
verify(op === 'b00100000, "Assert 857 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 858 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 859 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 216
#2;

verify(ir === 'b0000, "Assert 860 : < ir !== 'b0000 >");	// Vector No: 215
verify(op === 'b00000000, "Assert 861 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 862 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 863 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000000000000000000000000000000:0:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 217
#2;

verify(ir === 'b0000, "Assert 864 : < ir !== 'b0000 >");	// Vector No: 216
verify(op === 'b00000100, "Assert 865 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 866 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 867 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 218
#2;

verify(ir === 'b0000, "Assert 868 : < ir !== 'b0000 >");	// Vector No: 217
verify(op === 'b00000000, "Assert 869 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 870 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 871 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000000000000000000000000000000:1:0:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 219
#2;

verify(ir === 'b0000, "Assert 872 : < ir !== 'b0000 >");	// Vector No: 218
verify(op === 'b01000000, "Assert 873 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 874 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 875 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 220
#2;

verify(ir === 'b0000, "Assert 876 : < ir !== 'b0000 >");	// Vector No: 219
verify(op === 'b00000000, "Assert 877 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 878 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 879 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 221
#2;

verify(ir === 'b0000, "Assert 880 : < ir !== 'b0000 >");	// Vector No: 220
verify(op === 'b00001000, "Assert 881 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 882 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 883 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 222
#2;

verify(ir === 'b0000, "Assert 884 : < ir !== 'b0000 >");	// Vector No: 221
verify(op === 'b00000000, "Assert 885 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 886 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 887 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 223
#2;

verify(ir === 'b0000, "Assert 888 : < ir !== 'b0000 >");	// Vector No: 222
verify(op === 'b10000000, "Assert 889 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 890 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 891 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 224
#2;

verify(ir === 'b0000, "Assert 892 : < ir !== 'b0000 >");	// Vector No: 223
verify(op === 'b00000000, "Assert 893 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 894 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 895 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000000000000000000000000000000:0:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 225
#2;

verify(ir === 'b0000, "Assert 896 : < ir !== 'b0000 >");	// Vector No: 224
verify(op === 'b00010000, "Assert 897 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 898 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 899 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 226
#2;

verify(ir === 'b0000, "Assert 900 : < ir !== 'b0000 >");	// Vector No: 225
verify(op === 'b00000000, "Assert 901 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 902 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 903 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000000000000000000000000000000:1:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 227
#2;

verify(ir === 'b0001, "Assert 904 : < ir !== 'b0001 >");	// Vector No: 226
verify(op === 'b00000000, "Assert 905 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 906 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 907 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 228
#2;

verify(ir === 'b0000, "Assert 908 : < ir !== 'b0000 >");	// Vector No: 227
verify(op === 'b00000000, "Assert 909 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 910 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 911 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000000000000000000000000000000:0:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 229
#2;

verify(ir === 'b0000, "Assert 912 : < ir !== 'b0000 >");	// Vector No: 228
verify(op === 'b00100000, "Assert 913 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 914 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 915 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 230
#2;

verify(ir === 'b0000, "Assert 916 : < ir !== 'b0000 >");	// Vector No: 229
verify(op === 'b00000000, "Assert 917 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 918 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 919 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000000000000000000000000000000:1:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 231
#2;

verify(ir === 'b0010, "Assert 920 : < ir !== 'b0010 >");	// Vector No: 230
verify(op === 'b00000000, "Assert 921 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 922 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 923 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 232
#2;

verify(ir === 'b0000, "Assert 924 : < ir !== 'b0000 >");	// Vector No: 231
verify(op === 'b00000000, "Assert 925 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 926 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 927 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000000000000000000000000000000:0:0:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 233
#2;

verify(ir === 'b0000, "Assert 928 : < ir !== 'b0000 >");	// Vector No: 232
verify(op === 'b01000000, "Assert 929 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 930 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 931 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 234
#2;

verify(ir === 'b0000, "Assert 932 : < ir !== 'b0000 >");	// Vector No: 233
verify(op === 'b00000000, "Assert 933 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 934 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 935 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000000000000000000000000000000:1:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 235
#2;

verify(ir === 'b0100, "Assert 936 : < ir !== 'b0100 >");	// Vector No: 234
verify(op === 'b00000000, "Assert 937 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 938 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 939 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 236
#2;

verify(ir === 'b0000, "Assert 940 : < ir !== 'b0000 >");	// Vector No: 235
verify(op === 'b00000000, "Assert 941 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 942 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 943 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000000000000000000000000000000:0:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 237
#2;

verify(ir === 'b0000, "Assert 944 : < ir !== 'b0000 >");	// Vector No: 236
verify(op === 'b10000000, "Assert 945 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 946 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 947 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 238
#2;

verify(ir === 'b0000, "Assert 948 : < ir !== 'b0000 >");	// Vector No: 237
verify(op === 'b00000000, "Assert 949 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 950 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 951 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 239
#2;

verify(ir === 'b0000, "Assert 952 : < ir !== 'b0000 >");	// Vector No: 238
verify(op === 'b00000000, "Assert 953 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 954 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 955 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 240
#2;

verify(ir === 'b0000, "Assert 956 : < ir !== 'b0000 >");	// Vector No: 239
verify(op === 'b00000000, "Assert 957 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 958 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 959 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000000000000000000000000000000:0:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 241
#2;

verify(ir === 'b0001, "Assert 960 : < ir !== 'b0001 >");	// Vector No: 240
verify(op === 'b00000000, "Assert 961 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 962 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 963 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 242
#2;

verify(ir === 'b0000, "Assert 964 : < ir !== 'b0000 >");	// Vector No: 241
verify(op === 'b00000000, "Assert 965 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 966 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 967 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 243
#2;

verify(ir === 'b0000, "Assert 968 : < ir !== 'b0000 >");	// Vector No: 242
verify(op === 'b00000000, "Assert 969 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 970 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 971 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 244
#2;

verify(ir === 'b0000, "Assert 972 : < ir !== 'b0000 >");	// Vector No: 243
verify(op === 'b00000000, "Assert 973 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 974 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 975 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000000000000000000000000000000:0:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 245
#2;

verify(ir === 'b0010, "Assert 976 : < ir !== 'b0010 >");	// Vector No: 244
verify(op === 'b00000000, "Assert 977 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 978 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 979 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 246
#2;

verify(ir === 'b0000, "Assert 980 : < ir !== 'b0000 >");	// Vector No: 245
verify(op === 'b00000000, "Assert 981 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 982 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 983 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 247
#2;

verify(ir === 'b0000, "Assert 984 : < ir !== 'b0000 >");	// Vector No: 246
verify(op === 'b00000000, "Assert 985 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 986 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 987 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 248
#2;

verify(ir === 'b0000, "Assert 988 : < ir !== 'b0000 >");	// Vector No: 247
verify(op === 'b00000000, "Assert 989 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 990 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 991 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000000000000000000000000000000:0:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 249
#2;

verify(ir === 'b0100, "Assert 992 : < ir !== 'b0100 >");	// Vector No: 248
verify(op === 'b00000000, "Assert 993 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 994 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 995 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 250
#2;

verify(ir === 'b0000, "Assert 996 : < ir !== 'b0000 >");	// Vector No: 249
verify(op === 'b00000000, "Assert 997 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 998 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 999 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 251
#2;

verify(ir === 'b0000, "Assert 1000 : < ir !== 'b0000 >");	// Vector No: 250
verify(op === 'b00000000, "Assert 1001 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1002 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1003 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 252
#2;

verify(ir === 'b0000, "Assert 1004 : < ir !== 'b0000 >");	// Vector No: 251
verify(op === 'b00000000, "Assert 1005 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1006 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1007 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000000000000000000000000000000:0:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 253
#2;

verify(ir === 'b1000, "Assert 1008 : < ir !== 'b1000 >");	// Vector No: 252
verify(op === 'b00000000, "Assert 1009 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1010 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1011 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 254
#2;

verify(ir === 'b0000, "Assert 1012 : < ir !== 'b0000 >");	// Vector No: 253
verify(op === 'b00000000, "Assert 1013 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1014 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1015 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000000000000000000000000000000:1:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 255
#2;

verify(ir === 'b1000, "Assert 1016 : < ir !== 'b1000 >");	// Vector No: 254
verify(op === 'b00000000, "Assert 1017 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1018 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1019 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 256
#2;

verify(ir === 'b0000, "Assert 1020 : < ir !== 'b0000 >");	// Vector No: 255
verify(op === 'b00000000, "Assert 1021 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 1022 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 1023 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111110:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111110;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 257
#2;

verify(ir === 'b1111, "Assert 1024 : < ir !== 'b1111 >");	// Vector No: 256
verify(op === 'b11111111, "Assert 1025 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1026 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1027 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111110:0:1:1111:11111111:0:11111111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111110;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 258
#2;

verify(ir === 'b1111, "Assert 1028 : < ir !== 'b1111 >");	// Vector No: 257
verify(op === 'b11111111, "Assert 1029 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1030 : < extop !== 0 >");
verify(addr === 'b11111111111111111110, "Assert 1031 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111110:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111110;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 259
#2;

verify(ir === 'b1111, "Assert 1032 : < ir !== 'b1111 >");	// Vector No: 258
verify(op === 'b11111000, "Assert 1033 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1034 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1035 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111110:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111110;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 260
#2;

verify(ir === 'b1111, "Assert 1036 : < ir !== 'b1111 >");	// Vector No: 259
verify(op === 'b11111000, "Assert 1037 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1038 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1039 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111101:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111101;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 261
#2;

verify(ir === 'b1111, "Assert 1040 : < ir !== 'b1111 >");	// Vector No: 260
verify(op === 'b11111111, "Assert 1041 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1042 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1043 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111101:0:1:1111:11111111:0:11111111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111101;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 262
#2;

verify(ir === 'b1111, "Assert 1044 : < ir !== 'b1111 >");	// Vector No: 261
verify(op === 'b11111111, "Assert 1045 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1046 : < extop !== 0 >");
verify(addr === 'b11111111111111111101, "Assert 1047 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111101:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111101;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 263
#2;

verify(ir === 'b1111, "Assert 1048 : < ir !== 'b1111 >");	// Vector No: 262
verify(op === 'b11111000, "Assert 1049 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1050 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1051 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111101:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111101;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 264
#2;

verify(ir === 'b1111, "Assert 1052 : < ir !== 'b1111 >");	// Vector No: 263
verify(op === 'b11111000, "Assert 1053 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1054 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1055 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111011:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111011;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 265
#2;

verify(ir === 'b1111, "Assert 1056 : < ir !== 'b1111 >");	// Vector No: 264
verify(op === 'b11111111, "Assert 1057 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1058 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1059 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111011:0:1:1111:11111111:0:11111111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111011;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 266
#2;

verify(ir === 'b1111, "Assert 1060 : < ir !== 'b1111 >");	// Vector No: 265
verify(op === 'b11111111, "Assert 1061 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1062 : < extop !== 0 >");
verify(addr === 'b11111111111111111011, "Assert 1063 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111011:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111011;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 267
#2;

verify(ir === 'b1111, "Assert 1064 : < ir !== 'b1111 >");	// Vector No: 266
verify(op === 'b11111000, "Assert 1065 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1066 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1067 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111111011:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111111011;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 268
#2;

verify(ir === 'b1111, "Assert 1068 : < ir !== 'b1111 >");	// Vector No: 267
verify(op === 'b11111000, "Assert 1069 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1070 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1071 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111110111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111110111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 269
#2;

verify(ir === 'b1111, "Assert 1072 : < ir !== 'b1111 >");	// Vector No: 268
verify(op === 'b11111111, "Assert 1073 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1074 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1075 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111110111:0:1:1111:11111111:0:11111111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111110111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 270
#2;

verify(ir === 'b1111, "Assert 1076 : < ir !== 'b1111 >");	// Vector No: 269
verify(op === 'b11111111, "Assert 1077 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1078 : < extop !== 0 >");
verify(addr === 'b11111111111111110111, "Assert 1079 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111110111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111110111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 271
#2;

verify(ir === 'b1111, "Assert 1080 : < ir !== 'b1111 >");	// Vector No: 270
verify(op === 'b11111000, "Assert 1081 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1082 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1083 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111110111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111110111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 272
#2;

verify(ir === 'b1111, "Assert 1084 : < ir !== 'b1111 >");	// Vector No: 271
verify(op === 'b11111000, "Assert 1085 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1086 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1087 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111101111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111101111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 273
#2;

verify(ir === 'b1111, "Assert 1088 : < ir !== 'b1111 >");	// Vector No: 272
verify(op === 'b11111111, "Assert 1089 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1090 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1091 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111101111:0:1:1111:11111111:0:11111111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111101111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 274
#2;

verify(ir === 'b1111, "Assert 1092 : < ir !== 'b1111 >");	// Vector No: 273
verify(op === 'b11111111, "Assert 1093 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1094 : < extop !== 0 >");
verify(addr === 'b11111111111111101111, "Assert 1095 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111101111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111101111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 275
#2;

verify(ir === 'b1111, "Assert 1096 : < ir !== 'b1111 >");	// Vector No: 274
verify(op === 'b11111000, "Assert 1097 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1098 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1099 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111101111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111101111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 276
#2;

verify(ir === 'b1111, "Assert 1100 : < ir !== 'b1111 >");	// Vector No: 275
verify(op === 'b11111000, "Assert 1101 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1102 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1103 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111011111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111011111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 277
#2;

verify(ir === 'b1111, "Assert 1104 : < ir !== 'b1111 >");	// Vector No: 276
verify(op === 'b11111111, "Assert 1105 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1106 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1107 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111011111:0:1:1111:11111111:0:11111111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111011111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 278
#2;

verify(ir === 'b1111, "Assert 1108 : < ir !== 'b1111 >");	// Vector No: 277
verify(op === 'b11111111, "Assert 1109 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1110 : < extop !== 0 >");
verify(addr === 'b11111111111111011111, "Assert 1111 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111011111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111011111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 279
#2;

verify(ir === 'b1111, "Assert 1112 : < ir !== 'b1111 >");	// Vector No: 278
verify(op === 'b11111000, "Assert 1113 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1114 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1115 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111111011111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111111011111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 280
#2;

verify(ir === 'b1111, "Assert 1116 : < ir !== 'b1111 >");	// Vector No: 279
verify(op === 'b11111000, "Assert 1117 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1118 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1119 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111110111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111110111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 281
#2;

verify(ir === 'b1111, "Assert 1120 : < ir !== 'b1111 >");	// Vector No: 280
verify(op === 'b11111111, "Assert 1121 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1122 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1123 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111110111111:0:1:1111:11111111:0:11111111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111110111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 282
#2;

verify(ir === 'b1111, "Assert 1124 : < ir !== 'b1111 >");	// Vector No: 281
verify(op === 'b11111111, "Assert 1125 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1126 : < extop !== 0 >");
verify(addr === 'b11111111111110111111, "Assert 1127 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111110111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111110111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 283
#2;

verify(ir === 'b1111, "Assert 1128 : < ir !== 'b1111 >");	// Vector No: 282
verify(op === 'b11111000, "Assert 1129 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1130 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1131 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111110111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111110111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 284
#2;

verify(ir === 'b1111, "Assert 1132 : < ir !== 'b1111 >");	// Vector No: 283
verify(op === 'b11111000, "Assert 1133 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1134 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1135 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111101111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111101111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 285
#2;

verify(ir === 'b1111, "Assert 1136 : < ir !== 'b1111 >");	// Vector No: 284
verify(op === 'b11111111, "Assert 1137 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1138 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1139 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111101111111:0:1:1111:11111111:0:11111111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111101111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 286
#2;

verify(ir === 'b1111, "Assert 1140 : < ir !== 'b1111 >");	// Vector No: 285
verify(op === 'b11111111, "Assert 1141 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1142 : < extop !== 0 >");
verify(addr === 'b11111111111101111111, "Assert 1143 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111101111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111101111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 287
#2;

verify(ir === 'b1111, "Assert 1144 : < ir !== 'b1111 >");	// Vector No: 286
verify(op === 'b11111000, "Assert 1145 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1146 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1147 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111101111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111101111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 288
#2;

verify(ir === 'b1111, "Assert 1148 : < ir !== 'b1111 >");	// Vector No: 287
verify(op === 'b11111000, "Assert 1149 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1150 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1151 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111011111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111011111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 289
#2;

verify(ir === 'b1111, "Assert 1152 : < ir !== 'b1111 >");	// Vector No: 288
verify(op === 'b11111111, "Assert 1153 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1154 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1155 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111011111111:0:1:1111:11111111:0:11111111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111011111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 290
#2;

verify(ir === 'b1111, "Assert 1156 : < ir !== 'b1111 >");	// Vector No: 289
verify(op === 'b11111111, "Assert 1157 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1158 : < extop !== 0 >");
verify(addr === 'b11111111111011111111, "Assert 1159 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111011111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111011111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 291
#2;

verify(ir === 'b1111, "Assert 1160 : < ir !== 'b1111 >");	// Vector No: 290
verify(op === 'b11111000, "Assert 1161 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1162 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1163 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111111011111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111111011111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 292
#2;

verify(ir === 'b1111, "Assert 1164 : < ir !== 'b1111 >");	// Vector No: 291
verify(op === 'b11111000, "Assert 1165 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1166 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1167 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111110111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111110111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 293
#2;

verify(ir === 'b1111, "Assert 1168 : < ir !== 'b1111 >");	// Vector No: 292
verify(op === 'b11111111, "Assert 1169 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1170 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1171 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111110111111111:0:1:1111:11111111:0:11111111110111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111110111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 294
#2;

verify(ir === 'b1111, "Assert 1172 : < ir !== 'b1111 >");	// Vector No: 293
verify(op === 'b11111111, "Assert 1173 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1174 : < extop !== 0 >");
verify(addr === 'b11111111110111111111, "Assert 1175 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111110111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111110111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 295
#2;

verify(ir === 'b1111, "Assert 1176 : < ir !== 'b1111 >");	// Vector No: 294
verify(op === 'b11111000, "Assert 1177 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1178 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1179 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111110111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111110111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 296
#2;

verify(ir === 'b1111, "Assert 1180 : < ir !== 'b1111 >");	// Vector No: 295
verify(op === 'b11111000, "Assert 1181 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1182 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1183 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111101111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111101111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 297
#2;

verify(ir === 'b1111, "Assert 1184 : < ir !== 'b1111 >");	// Vector No: 296
verify(op === 'b11111111, "Assert 1185 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1186 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1187 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111101111111111:0:1:1111:11111111:0:11111111101111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111101111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 298
#2;

verify(ir === 'b1111, "Assert 1188 : < ir !== 'b1111 >");	// Vector No: 297
verify(op === 'b11111111, "Assert 1189 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1190 : < extop !== 0 >");
verify(addr === 'b11111111101111111111, "Assert 1191 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111101111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111101111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 299
#2;

verify(ir === 'b1111, "Assert 1192 : < ir !== 'b1111 >");	// Vector No: 298
verify(op === 'b11111000, "Assert 1193 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1194 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1195 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111101111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111101111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 300
#2;

verify(ir === 'b1111, "Assert 1196 : < ir !== 'b1111 >");	// Vector No: 299
verify(op === 'b11111000, "Assert 1197 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1198 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1199 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111011111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111011111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 301
#2;

verify(ir === 'b1111, "Assert 1200 : < ir !== 'b1111 >");	// Vector No: 300
verify(op === 'b11111111, "Assert 1201 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1202 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1203 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111011111111111:0:1:1111:11111111:0:11111111011111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111011111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 302
#2;

verify(ir === 'b1111, "Assert 1204 : < ir !== 'b1111 >");	// Vector No: 301
verify(op === 'b11111111, "Assert 1205 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1206 : < extop !== 0 >");
verify(addr === 'b11111111011111111111, "Assert 1207 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111011111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111011111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 303
#2;

verify(ir === 'b1111, "Assert 1208 : < ir !== 'b1111 >");	// Vector No: 302
verify(op === 'b11111000, "Assert 1209 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1210 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1211 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111111011111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111111011111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 304
#2;

verify(ir === 'b1111, "Assert 1212 : < ir !== 'b1111 >");	// Vector No: 303
verify(op === 'b11111000, "Assert 1213 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1214 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1215 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111110111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111110111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 305
#2;

verify(ir === 'b1111, "Assert 1216 : < ir !== 'b1111 >");	// Vector No: 304
verify(op === 'b11111111, "Assert 1217 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1218 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1219 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111110111111111111:0:1:1111:11111111:0:11111110111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111110111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 306
#2;

verify(ir === 'b1111, "Assert 1220 : < ir !== 'b1111 >");	// Vector No: 305
verify(op === 'b11111111, "Assert 1221 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1222 : < extop !== 0 >");
verify(addr === 'b11111110111111111111, "Assert 1223 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111110111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111110111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 307
#2;

verify(ir === 'b1111, "Assert 1224 : < ir !== 'b1111 >");	// Vector No: 306
verify(op === 'b11111000, "Assert 1225 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1226 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1227 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111110111111111111:1:1:1111:11111000:0:00000111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111110111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 308
#2;

verify(ir === 'b1111, "Assert 1228 : < ir !== 'b1111 >");	// Vector No: 307
verify(op === 'b11111000, "Assert 1229 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1230 : < extop !== 0 >");
verify(addr === 'b00000111111111111110, "Assert 1231 : < addr !== 'b00000111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111101111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111101111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 309
#2;

verify(ir === 'b1111, "Assert 1232 : < ir !== 'b1111 >");	// Vector No: 308
verify(op === 'b11111111, "Assert 1233 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1234 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1235 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111101111111111111:0:1:1111:11111111:0:11111101111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111101111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 310
#2;

verify(ir === 'b1111, "Assert 1236 : < ir !== 'b1111 >");	// Vector No: 309
verify(op === 'b11111111, "Assert 1237 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1238 : < extop !== 0 >");
verify(addr === 'b11111101111111111111, "Assert 1239 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111101111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111101111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 311
#2;

verify(ir === 'b1111, "Assert 1240 : < ir !== 'b1111 >");	// Vector No: 310
verify(op === 'b11111000, "Assert 1241 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1242 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1243 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111101111111111111:1:1:1111:11111000:0:00000111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111101111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 312
#2;

verify(ir === 'b1111, "Assert 1244 : < ir !== 'b1111 >");	// Vector No: 311
verify(op === 'b11111000, "Assert 1245 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1246 : < extop !== 0 >");
verify(addr === 'b00000111111111111101, "Assert 1247 : < addr !== 'b00000111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111011111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111011111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 313
#2;

verify(ir === 'b1111, "Assert 1248 : < ir !== 'b1111 >");	// Vector No: 312
verify(op === 'b11111111, "Assert 1249 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1250 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1251 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111011111111111111:0:1:1111:11111111:0:11111011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111011111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 314
#2;

verify(ir === 'b1111, "Assert 1252 : < ir !== 'b1111 >");	// Vector No: 313
verify(op === 'b11111111, "Assert 1253 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1254 : < extop !== 0 >");
verify(addr === 'b11111011111111111111, "Assert 1255 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111011111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111011111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 315
#2;

verify(ir === 'b1111, "Assert 1256 : < ir !== 'b1111 >");	// Vector No: 314
verify(op === 'b11111000, "Assert 1257 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1258 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1259 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111111011111111111111:1:1:1111:11111000:0:00000111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111111011111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 316
#2;

verify(ir === 'b1111, "Assert 1260 : < ir !== 'b1111 >");	// Vector No: 315
verify(op === 'b11111000, "Assert 1261 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1262 : < extop !== 0 >");
verify(addr === 'b00000111111111111011, "Assert 1263 : < addr !== 'b00000111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111110111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111110111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 317
#2;

verify(ir === 'b1111, "Assert 1264 : < ir !== 'b1111 >");	// Vector No: 316
verify(op === 'b11111111, "Assert 1265 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1266 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1267 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111110111111111111111:0:1:1111:11111111:0:11110111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111110111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 318
#2;

verify(ir === 'b1111, "Assert 1268 : < ir !== 'b1111 >");	// Vector No: 317
verify(op === 'b11111111, "Assert 1269 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1270 : < extop !== 0 >");
verify(addr === 'b11110111111111111111, "Assert 1271 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111110111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111110111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 319
#2;

verify(ir === 'b1111, "Assert 1272 : < ir !== 'b1111 >");	// Vector No: 318
verify(op === 'b11111000, "Assert 1273 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1274 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1275 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111110111111111111111:1:1:1111:11111000:0:00000111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111110111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 320
#2;

verify(ir === 'b1111, "Assert 1276 : < ir !== 'b1111 >");	// Vector No: 319
verify(op === 'b11111000, "Assert 1277 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1278 : < extop !== 0 >");
verify(addr === 'b00000111111111110111, "Assert 1279 : < addr !== 'b00000111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111101111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111101111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 321
#2;

verify(ir === 'b1111, "Assert 1280 : < ir !== 'b1111 >");	// Vector No: 320
verify(op === 'b11111111, "Assert 1281 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1282 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1283 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111101111111111111111:0:1:1111:11111111:0:11101111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111101111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 322
#2;

verify(ir === 'b1111, "Assert 1284 : < ir !== 'b1111 >");	// Vector No: 321
verify(op === 'b11111111, "Assert 1285 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1286 : < extop !== 0 >");
verify(addr === 'b11101111111111111111, "Assert 1287 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111101111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111101111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 323
#2;

verify(ir === 'b1111, "Assert 1288 : < ir !== 'b1111 >");	// Vector No: 322
verify(op === 'b11111000, "Assert 1289 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1290 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1291 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111101111111111111111:1:1:1111:11111000:0:00000111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111101111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 324
#2;

verify(ir === 'b1111, "Assert 1292 : < ir !== 'b1111 >");	// Vector No: 323
verify(op === 'b11111000, "Assert 1293 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1294 : < extop !== 0 >");
verify(addr === 'b00000111111111101111, "Assert 1295 : < addr !== 'b00000111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111011111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111011111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 325
#2;

verify(ir === 'b1111, "Assert 1296 : < ir !== 'b1111 >");	// Vector No: 324
verify(op === 'b11111111, "Assert 1297 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1298 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1299 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111011111111111111111:0:1:1111:11111111:0:11011111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111011111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 326
#2;

verify(ir === 'b1111, "Assert 1300 : < ir !== 'b1111 >");	// Vector No: 325
verify(op === 'b11111111, "Assert 1301 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1302 : < extop !== 0 >");
verify(addr === 'b11011111111111111111, "Assert 1303 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111011111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111011111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 327
#2;

verify(ir === 'b1111, "Assert 1304 : < ir !== 'b1111 >");	// Vector No: 326
verify(op === 'b11111000, "Assert 1305 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1306 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1307 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111111011111111111111111:1:1:1111:11111000:0:00000111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111111011111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 328
#2;

verify(ir === 'b1111, "Assert 1308 : < ir !== 'b1111 >");	// Vector No: 327
verify(op === 'b11111000, "Assert 1309 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1310 : < extop !== 0 >");
verify(addr === 'b00000111111111011111, "Assert 1311 : < addr !== 'b00000111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111110111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111110111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 329
#2;

verify(ir === 'b1111, "Assert 1312 : < ir !== 'b1111 >");	// Vector No: 328
verify(op === 'b11111111, "Assert 1313 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1314 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1315 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111110111111111111111111:0:1:1111:11111111:0:10111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111110111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 330
#2;

verify(ir === 'b1111, "Assert 1316 : < ir !== 'b1111 >");	// Vector No: 329
verify(op === 'b11111111, "Assert 1317 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1318 : < extop !== 0 >");
verify(addr === 'b10111111111111111111, "Assert 1319 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111110111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111110111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 331
#2;

verify(ir === 'b1111, "Assert 1320 : < ir !== 'b1111 >");	// Vector No: 330
verify(op === 'b11111000, "Assert 1321 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1322 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1323 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111110111111111111111111:1:1:1111:11111000:0:00000111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111110111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 332
#2;

verify(ir === 'b1111, "Assert 1324 : < ir !== 'b1111 >");	// Vector No: 331
verify(op === 'b11111000, "Assert 1325 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1326 : < extop !== 0 >");
verify(addr === 'b00000111111110111111, "Assert 1327 : < addr !== 'b00000111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111101111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111101111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 333
#2;

verify(ir === 'b1111, "Assert 1328 : < ir !== 'b1111 >");	// Vector No: 332
verify(op === 'b11111111, "Assert 1329 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1330 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1331 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111101111111111111111111:0:1:1111:11111111:0:01111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111101111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 334
#2;

verify(ir === 'b1111, "Assert 1332 : < ir !== 'b1111 >");	// Vector No: 333
verify(op === 'b11111111, "Assert 1333 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1334 : < extop !== 0 >");
verify(addr === 'b01111111111111111111, "Assert 1335 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111101111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111101111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 335
#2;

verify(ir === 'b1111, "Assert 1336 : < ir !== 'b1111 >");	// Vector No: 334
verify(op === 'b11111000, "Assert 1337 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1338 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1339 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111101111111111111111111:1:1:1111:11111000:0:00000111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111101111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 336
#2;

verify(ir === 'b1111, "Assert 1340 : < ir !== 'b1111 >");	// Vector No: 335
verify(op === 'b11111000, "Assert 1341 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1342 : < extop !== 0 >");
verify(addr === 'b00000111111101111111, "Assert 1343 : < addr !== 'b00000111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111011111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111011111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 337
#2;

verify(ir === 'b1111, "Assert 1344 : < ir !== 'b1111 >");	// Vector No: 336
verify(op === 'b11111111, "Assert 1345 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1346 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1347 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111011111111111111111111:0:1:1111:11111110:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111011111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 338
#2;

verify(ir === 'b1111, "Assert 1348 : < ir !== 'b1111 >");	// Vector No: 337
verify(op === 'b11111110, "Assert 1349 : < op !== 'b11111110 >");
verify(extop === 0, "Assert 1350 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1351 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111011111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111011111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 339
#2;

verify(ir === 'b1111, "Assert 1352 : < ir !== 'b1111 >");	// Vector No: 338
verify(op === 'b11111000, "Assert 1353 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1354 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1355 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111111011111111111111111111:1:1:1111:11111000:0:00000111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111111011111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 340
#2;

verify(ir === 'b1111, "Assert 1356 : < ir !== 'b1111 >");	// Vector No: 339
verify(op === 'b11111000, "Assert 1357 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1358 : < extop !== 0 >");
verify(addr === 'b00000111111011111111, "Assert 1359 : < addr !== 'b00000111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111110111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111110111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 341
#2;

verify(ir === 'b1111, "Assert 1360 : < ir !== 'b1111 >");	// Vector No: 340
verify(op === 'b11111111, "Assert 1361 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1362 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1363 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111110111111111111111111111:0:1:1111:11111101:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111110111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 342
#2;

verify(ir === 'b1111, "Assert 1364 : < ir !== 'b1111 >");	// Vector No: 341
verify(op === 'b11111101, "Assert 1365 : < op !== 'b11111101 >");
verify(extop === 0, "Assert 1366 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1367 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111110111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111110111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 343
#2;

verify(ir === 'b1111, "Assert 1368 : < ir !== 'b1111 >");	// Vector No: 342
verify(op === 'b11111000, "Assert 1369 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1370 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1371 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111110111111111111111111111:1:1:1111:11111000:0:00000111110111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111110111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 344
#2;

verify(ir === 'b1111, "Assert 1372 : < ir !== 'b1111 >");	// Vector No: 343
verify(op === 'b11111000, "Assert 1373 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1374 : < extop !== 0 >");
verify(addr === 'b00000111110111111111, "Assert 1375 : < addr !== 'b00000111110111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111101111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111101111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 345
#2;

verify(ir === 'b1111, "Assert 1376 : < ir !== 'b1111 >");	// Vector No: 344
verify(op === 'b11111111, "Assert 1377 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1378 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1379 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111101111111111111111111111:0:1:1111:11111011:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111101111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 346
#2;

verify(ir === 'b1111, "Assert 1380 : < ir !== 'b1111 >");	// Vector No: 345
verify(op === 'b11111011, "Assert 1381 : < op !== 'b11111011 >");
verify(extop === 0, "Assert 1382 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1383 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111101111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111101111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 347
#2;

verify(ir === 'b1111, "Assert 1384 : < ir !== 'b1111 >");	// Vector No: 346
verify(op === 'b11111000, "Assert 1385 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1386 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1387 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111101111111111111111111111:1:1:1111:11111000:0:00000111101111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111101111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 348
#2;

verify(ir === 'b1111, "Assert 1388 : < ir !== 'b1111 >");	// Vector No: 347
verify(op === 'b11111000, "Assert 1389 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1390 : < extop !== 0 >");
verify(addr === 'b00000111101111111111, "Assert 1391 : < addr !== 'b00000111101111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111011111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111011111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 349
#2;

verify(ir === 'b1111, "Assert 1392 : < ir !== 'b1111 >");	// Vector No: 348
verify(op === 'b11111111, "Assert 1393 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1394 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1395 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111011111111111111111111111:0:1:1111:11110111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111011111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 350
#2;

verify(ir === 'b1111, "Assert 1396 : < ir !== 'b1111 >");	// Vector No: 349
verify(op === 'b11110111, "Assert 1397 : < op !== 'b11110111 >");
verify(extop === 0, "Assert 1398 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1399 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111011111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111011111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 351
#2;

verify(ir === 'b1111, "Assert 1400 : < ir !== 'b1111 >");	// Vector No: 350
verify(op === 'b11111000, "Assert 1401 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1402 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1403 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111111011111111111111111111111:1:1:1111:11111000:0:00000111011111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111111011111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 352
#2;

verify(ir === 'b1111, "Assert 1404 : < ir !== 'b1111 >");	// Vector No: 351
verify(op === 'b11111000, "Assert 1405 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1406 : < extop !== 0 >");
verify(addr === 'b00000111011111111111, "Assert 1407 : < addr !== 'b00000111011111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111110111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111110111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 353
#2;

verify(ir === 'b1111, "Assert 1408 : < ir !== 'b1111 >");	// Vector No: 352
verify(op === 'b11111111, "Assert 1409 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1410 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1411 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111110111111111111111111111111:0:1:1111:11101111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111110111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 354
#2;

verify(ir === 'b1111, "Assert 1412 : < ir !== 'b1111 >");	// Vector No: 353
verify(op === 'b11101111, "Assert 1413 : < op !== 'b11101111 >");
verify(extop === 0, "Assert 1414 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1415 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111110111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111110111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 355
#2;

verify(ir === 'b1111, "Assert 1416 : < ir !== 'b1111 >");	// Vector No: 354
verify(op === 'b11111000, "Assert 1417 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1418 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1419 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111110111111111111111111111111:1:1:1111:11111000:0:00000110111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111110111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 356
#2;

verify(ir === 'b1111, "Assert 1420 : < ir !== 'b1111 >");	// Vector No: 355
verify(op === 'b11111000, "Assert 1421 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1422 : < extop !== 0 >");
verify(addr === 'b00000110111111111111, "Assert 1423 : < addr !== 'b00000110111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111101111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111101111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 357
#2;

verify(ir === 'b1111, "Assert 1424 : < ir !== 'b1111 >");	// Vector No: 356
verify(op === 'b11111111, "Assert 1425 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1426 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1427 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111101111111111111111111111111:0:1:1111:11011111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111101111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 358
#2;

verify(ir === 'b1111, "Assert 1428 : < ir !== 'b1111 >");	// Vector No: 357
verify(op === 'b11011111, "Assert 1429 : < op !== 'b11011111 >");
verify(extop === 0, "Assert 1430 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1431 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111101111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111101111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 359
#2;

verify(ir === 'b1111, "Assert 1432 : < ir !== 'b1111 >");	// Vector No: 358
verify(op === 'b11111000, "Assert 1433 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1434 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1435 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111101111111111111111111111111:1:1:1111:11111000:0:00000101111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111101111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 360
#2;

verify(ir === 'b1111, "Assert 1436 : < ir !== 'b1111 >");	// Vector No: 359
verify(op === 'b11111000, "Assert 1437 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1438 : < extop !== 0 >");
verify(addr === 'b00000101111111111111, "Assert 1439 : < addr !== 'b00000101111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 361
#2;

verify(ir === 'b1111, "Assert 1440 : < ir !== 'b1111 >");	// Vector No: 360
verify(op === 'b11111111, "Assert 1441 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1442 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1443 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111011111111111111111111111111:0:1:1111:10111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 362
#2;

verify(ir === 'b1111, "Assert 1444 : < ir !== 'b1111 >");	// Vector No: 361
verify(op === 'b10111111, "Assert 1445 : < op !== 'b10111111 >");
verify(extop === 0, "Assert 1446 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1447 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 363
#2;

verify(ir === 'b1111, "Assert 1448 : < ir !== 'b1111 >");	// Vector No: 362
verify(op === 'b11111000, "Assert 1449 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1450 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1451 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111111011111111111111111111111111:1:1:1111:11110000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111111011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 364
#2;

verify(ir === 'b1111, "Assert 1452 : < ir !== 'b1111 >");	// Vector No: 363
verify(op === 'b11110000, "Assert 1453 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 1454 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 1455 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110111111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 365
#2;

verify(ir === 'b1111, "Assert 1456 : < ir !== 'b1111 >");	// Vector No: 364
verify(op === 'b11111111, "Assert 1457 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1458 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1459 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110111111111111111111111111111:0:1:1111:01111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 366
#2;

verify(ir === 'b1111, "Assert 1460 : < ir !== 'b1111 >");	// Vector No: 365
verify(op === 'b01111111, "Assert 1461 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 1462 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1463 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 367
#2;

verify(ir === 'b1111, "Assert 1464 : < ir !== 'b1111 >");	// Vector No: 366
verify(op === 'b11111000, "Assert 1465 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1466 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1467 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110111111111111111111111111111:1:1:1111:11101000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 368
#2;

verify(ir === 'b1111, "Assert 1468 : < ir !== 'b1111 >");	// Vector No: 367
verify(op === 'b11101000, "Assert 1469 : < op !== 'b11101000 >");
verify(extop === 0, "Assert 1470 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1471 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111101111111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111101111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 369
#2;

verify(ir === 'b1111, "Assert 1472 : < ir !== 'b1111 >");	// Vector No: 368
verify(op === 'b11111111, "Assert 1473 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1474 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1475 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111101111111111111111111111111111:0:1:1110:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111101111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 370
#2;

verify(ir === 'b1110, "Assert 1476 : < ir !== 'b1110 >");	// Vector No: 369
verify(op === 'b11111111, "Assert 1477 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1478 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1479 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111101111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111101111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 371
#2;

verify(ir === 'b1111, "Assert 1480 : < ir !== 'b1111 >");	// Vector No: 370
verify(op === 'b11111000, "Assert 1481 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1482 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1483 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111101111111111111111111111111111:1:1:1111:11011000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111101111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 372
#2;

verify(ir === 'b1111, "Assert 1484 : < ir !== 'b1111 >");	// Vector No: 371
verify(op === 'b11011000, "Assert 1485 : < op !== 'b11011000 >");
verify(extop === 0, "Assert 1486 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1487 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111011111111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111011111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 373
#2;

verify(ir === 'b1111, "Assert 1488 : < ir !== 'b1111 >");	// Vector No: 372
verify(op === 'b11111111, "Assert 1489 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1490 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1491 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111011111111111111111111111111111:0:1:1101:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111011111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 374
#2;

verify(ir === 'b1101, "Assert 1492 : < ir !== 'b1101 >");	// Vector No: 373
verify(op === 'b11111111, "Assert 1493 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1494 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1495 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111011111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111011111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 375
#2;

verify(ir === 'b1111, "Assert 1496 : < ir !== 'b1111 >");	// Vector No: 374
verify(op === 'b11111000, "Assert 1497 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1498 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1499 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111011111111111111111111111111111:1:1:1111:10111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111011111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 376
#2;

verify(ir === 'b1111, "Assert 1500 : < ir !== 'b1111 >");	// Vector No: 375
verify(op === 'b10111000, "Assert 1501 : < op !== 'b10111000 >");
verify(extop === 0, "Assert 1502 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1503 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110111111111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 377
#2;

verify(ir === 'b1111, "Assert 1504 : < ir !== 'b1111 >");	// Vector No: 376
verify(op === 'b11111111, "Assert 1505 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1506 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1507 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110111111111111111111111111111111:0:1:1011:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 378
#2;

verify(ir === 'b1011, "Assert 1508 : < ir !== 'b1011 >");	// Vector No: 377
verify(op === 'b11111111, "Assert 1509 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1510 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1511 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 379
#2;

verify(ir === 'b1111, "Assert 1512 : < ir !== 'b1111 >");	// Vector No: 378
verify(op === 'b11111000, "Assert 1513 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1514 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1515 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110111111111111111111111111111111:1:1:1111:01111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 380
#2;

verify(ir === 'b1111, "Assert 1516 : < ir !== 'b1111 >");	// Vector No: 379
verify(op === 'b01111000, "Assert 1517 : < op !== 'b01111000 >");
verify(extop === 0, "Assert 1518 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1519 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101111111111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 381
#2;

verify(ir === 'b1111, "Assert 1520 : < ir !== 'b1111 >");	// Vector No: 380
verify(op === 'b11111111, "Assert 1521 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1522 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1523 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101111111111111111111111111111111:0:1:0111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 382
#2;

verify(ir === 'b0111, "Assert 1524 : < ir !== 'b0111 >");	// Vector No: 381
verify(op === 'b11111111, "Assert 1525 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1526 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1527 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 383
#2;

verify(ir === 'b1111, "Assert 1528 : < ir !== 'b1111 >");	// Vector No: 382
verify(op === 'b11111000, "Assert 1529 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1530 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1531 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101111111111111111111111111111111:1:1:1111:01111111:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 384
#2;

verify(ir === 'b1111, "Assert 1532 : < ir !== 'b1111 >");	// Vector No: 383
verify(op === 'b01111111, "Assert 1533 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 1534 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1535 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011111111111111111111111111111111:0:0:1111:11111111:0:11111111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 385
#2;

verify(ir === 'b1111, "Assert 1536 : < ir !== 'b1111 >");	// Vector No: 384
verify(op === 'b11111111, "Assert 1537 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1538 : < extop !== 0 >");
verify(addr === 'b11111111111111111110, "Assert 1539 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 386
#2;

verify(ir === 'b1111, "Assert 1540 : < ir !== 'b1111 >");	// Vector No: 385
verify(op === 'b11111111, "Assert 1541 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1542 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1543 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 387
#2;

verify(ir === 'b1111, "Assert 1544 : < ir !== 'b1111 >");	// Vector No: 386
verify(op === 'b11111000, "Assert 1545 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1546 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1547 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011111111111111111111111111111111:1:1:1110:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 388
#2;

verify(ir === 'b1110, "Assert 1548 : < ir !== 'b1110 >");	// Vector No: 387
verify(op === 'b11111000, "Assert 1549 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1550 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1551 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111111111111111111111111111111111:0:0:1111:11111111:0:11111111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 389
#2;

verify(ir === 'b1111, "Assert 1552 : < ir !== 'b1111 >");	// Vector No: 388
verify(op === 'b11111111, "Assert 1553 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1554 : < extop !== 0 >");
verify(addr === 'b11111111111111111101, "Assert 1555 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 390
#2;

verify(ir === 'b1111, "Assert 1556 : < ir !== 'b1111 >");	// Vector No: 389
verify(op === 'b11111111, "Assert 1557 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1558 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1559 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 391
#2;

verify(ir === 'b1111, "Assert 1560 : < ir !== 'b1111 >");	// Vector No: 390
verify(op === 'b11111000, "Assert 1561 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1562 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1563 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111111111111111111111111111111111:1:1:1101:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 392
#2;

verify(ir === 'b1101, "Assert 1564 : < ir !== 'b1101 >");	// Vector No: 391
verify(op === 'b11111000, "Assert 1565 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1566 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1567 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111111111111111111111111111111111:0:0:1111:11111111:0:11111111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 393
#2;

verify(ir === 'b1111, "Assert 1568 : < ir !== 'b1111 >");	// Vector No: 392
verify(op === 'b11111111, "Assert 1569 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1570 : < extop !== 0 >");
verify(addr === 'b11111111111111111011, "Assert 1571 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 394
#2;

verify(ir === 'b1111, "Assert 1572 : < ir !== 'b1111 >");	// Vector No: 393
verify(op === 'b11111111, "Assert 1573 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1574 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1575 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 395
#2;

verify(ir === 'b1111, "Assert 1576 : < ir !== 'b1111 >");	// Vector No: 394
verify(op === 'b11111000, "Assert 1577 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1578 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1579 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111111111111111111111111111111111:1:1:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 396
#2;

verify(ir === 'b1011, "Assert 1580 : < ir !== 'b1011 >");	// Vector No: 395
verify(op === 'b11111000, "Assert 1581 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1582 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1583 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111111111111111111111111111111111:0:0:1111:11111111:0:11111111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 397
#2;

verify(ir === 'b1111, "Assert 1584 : < ir !== 'b1111 >");	// Vector No: 396
verify(op === 'b11111111, "Assert 1585 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1586 : < extop !== 0 >");
verify(addr === 'b11111111111111110111, "Assert 1587 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 398
#2;

verify(ir === 'b1111, "Assert 1588 : < ir !== 'b1111 >");	// Vector No: 397
verify(op === 'b11111111, "Assert 1589 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1590 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1591 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 399
#2;

verify(ir === 'b1111, "Assert 1592 : < ir !== 'b1111 >");	// Vector No: 398
verify(op === 'b11111000, "Assert 1593 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1594 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1595 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111111111111111111111111111111111:1:1:0111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 400
#2;

verify(ir === 'b0111, "Assert 1596 : < ir !== 'b0111 >");	// Vector No: 399
verify(op === 'b11111000, "Assert 1597 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1598 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1599 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111111111111111111111111111111111:0:0:1111:11111111:0:11111111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 401
#2;

verify(ir === 'b1111, "Assert 1600 : < ir !== 'b1111 >");	// Vector No: 400
verify(op === 'b11111111, "Assert 1601 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1602 : < extop !== 0 >");
verify(addr === 'b11111111111111101111, "Assert 1603 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 402
#2;

verify(ir === 'b1111, "Assert 1604 : < ir !== 'b1111 >");	// Vector No: 401
verify(op === 'b11111111, "Assert 1605 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1606 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1607 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 403
#2;

verify(ir === 'b1111, "Assert 1608 : < ir !== 'b1111 >");	// Vector No: 402
verify(op === 'b11111000, "Assert 1609 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1610 : < extop !== 0 >");
verify(addr === 'b00000111111111111110, "Assert 1611 : < addr !== 'b00000111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 404
#2;

verify(ir === 'b1111, "Assert 1612 : < ir !== 'b1111 >");	// Vector No: 403
verify(op === 'b11111000, "Assert 1613 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1614 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1615 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111111111111111111111111111111111:0:0:1111:11111111:0:11111111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 405
#2;

verify(ir === 'b1111, "Assert 1616 : < ir !== 'b1111 >");	// Vector No: 404
verify(op === 'b11111111, "Assert 1617 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1618 : < extop !== 0 >");
verify(addr === 'b11111111111111011111, "Assert 1619 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 406
#2;

verify(ir === 'b1111, "Assert 1620 : < ir !== 'b1111 >");	// Vector No: 405
verify(op === 'b11111111, "Assert 1621 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1622 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1623 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 407
#2;

verify(ir === 'b1111, "Assert 1624 : < ir !== 'b1111 >");	// Vector No: 406
verify(op === 'b11111000, "Assert 1625 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1626 : < extop !== 0 >");
verify(addr === 'b00000111111111111101, "Assert 1627 : < addr !== 'b00000111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 408
#2;

verify(ir === 'b1111, "Assert 1628 : < ir !== 'b1111 >");	// Vector No: 407
verify(op === 'b11111000, "Assert 1629 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1630 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1631 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111111111111111111111111111111111:0:0:1111:11111111:0:11111111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 409
#2;

verify(ir === 'b1111, "Assert 1632 : < ir !== 'b1111 >");	// Vector No: 408
verify(op === 'b11111111, "Assert 1633 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1634 : < extop !== 0 >");
verify(addr === 'b11111111111110111111, "Assert 1635 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 410
#2;

verify(ir === 'b1111, "Assert 1636 : < ir !== 'b1111 >");	// Vector No: 409
verify(op === 'b11111111, "Assert 1637 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1638 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1639 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 411
#2;

verify(ir === 'b1111, "Assert 1640 : < ir !== 'b1111 >");	// Vector No: 410
verify(op === 'b11111000, "Assert 1641 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1642 : < extop !== 0 >");
verify(addr === 'b00000111111111111011, "Assert 1643 : < addr !== 'b00000111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 412
#2;

verify(ir === 'b1111, "Assert 1644 : < ir !== 'b1111 >");	// Vector No: 411
verify(op === 'b11111000, "Assert 1645 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1646 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1647 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111111111111111111111111111111111:0:0:1111:11111111:0:11111111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 413
#2;

verify(ir === 'b1111, "Assert 1648 : < ir !== 'b1111 >");	// Vector No: 412
verify(op === 'b11111111, "Assert 1649 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1650 : < extop !== 0 >");
verify(addr === 'b11111111111101111111, "Assert 1651 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 414
#2;

verify(ir === 'b1111, "Assert 1652 : < ir !== 'b1111 >");	// Vector No: 413
verify(op === 'b11111111, "Assert 1653 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1654 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1655 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 415
#2;

verify(ir === 'b1111, "Assert 1656 : < ir !== 'b1111 >");	// Vector No: 414
verify(op === 'b11111000, "Assert 1657 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1658 : < extop !== 0 >");
verify(addr === 'b00000111111111110111, "Assert 1659 : < addr !== 'b00000111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 416
#2;

verify(ir === 'b1111, "Assert 1660 : < ir !== 'b1111 >");	// Vector No: 415
verify(op === 'b11111000, "Assert 1661 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1662 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1663 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111111111111111111111111111111111:0:0:1111:11111111:0:11111111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 417
#2;

verify(ir === 'b1111, "Assert 1664 : < ir !== 'b1111 >");	// Vector No: 416
verify(op === 'b11111111, "Assert 1665 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1666 : < extop !== 0 >");
verify(addr === 'b11111111111011111111, "Assert 1667 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 418
#2;

verify(ir === 'b1111, "Assert 1668 : < ir !== 'b1111 >");	// Vector No: 417
verify(op === 'b11111111, "Assert 1669 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1670 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1671 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 419
#2;

verify(ir === 'b1111, "Assert 1672 : < ir !== 'b1111 >");	// Vector No: 418
verify(op === 'b11111000, "Assert 1673 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1674 : < extop !== 0 >");
verify(addr === 'b00000111111111101111, "Assert 1675 : < addr !== 'b00000111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 420
#2;

verify(ir === 'b1111, "Assert 1676 : < ir !== 'b1111 >");	// Vector No: 419
verify(op === 'b11111000, "Assert 1677 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1678 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1679 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111111111111111111111111111111111:0:0:1111:11111111:0:11111111110111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 421
#2;

verify(ir === 'b1111, "Assert 1680 : < ir !== 'b1111 >");	// Vector No: 420
verify(op === 'b11111111, "Assert 1681 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1682 : < extop !== 0 >");
verify(addr === 'b11111111110111111111, "Assert 1683 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 422
#2;

verify(ir === 'b1111, "Assert 1684 : < ir !== 'b1111 >");	// Vector No: 421
verify(op === 'b11111111, "Assert 1685 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1686 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1687 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 423
#2;

verify(ir === 'b1111, "Assert 1688 : < ir !== 'b1111 >");	// Vector No: 422
verify(op === 'b11111000, "Assert 1689 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1690 : < extop !== 0 >");
verify(addr === 'b00000111111111011111, "Assert 1691 : < addr !== 'b00000111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 424
#2;

verify(ir === 'b1111, "Assert 1692 : < ir !== 'b1111 >");	// Vector No: 423
verify(op === 'b11111000, "Assert 1693 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1694 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1695 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111111111111111111111111111111111:0:0:1111:11111111:0:11111111101111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 425
#2;

verify(ir === 'b1111, "Assert 1696 : < ir !== 'b1111 >");	// Vector No: 424
verify(op === 'b11111111, "Assert 1697 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1698 : < extop !== 0 >");
verify(addr === 'b11111111101111111111, "Assert 1699 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 426
#2;

verify(ir === 'b1111, "Assert 1700 : < ir !== 'b1111 >");	// Vector No: 425
verify(op === 'b11111111, "Assert 1701 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1702 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1703 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 427
#2;

verify(ir === 'b1111, "Assert 1704 : < ir !== 'b1111 >");	// Vector No: 426
verify(op === 'b11111000, "Assert 1705 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1706 : < extop !== 0 >");
verify(addr === 'b00000111111110111111, "Assert 1707 : < addr !== 'b00000111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 428
#2;

verify(ir === 'b1111, "Assert 1708 : < ir !== 'b1111 >");	// Vector No: 427
verify(op === 'b11111000, "Assert 1709 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1710 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1711 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111111111111111111111111111111111:0:0:1111:11111111:0:11111111011111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 429
#2;

verify(ir === 'b1111, "Assert 1712 : < ir !== 'b1111 >");	// Vector No: 428
verify(op === 'b11111111, "Assert 1713 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1714 : < extop !== 0 >");
verify(addr === 'b11111111011111111111, "Assert 1715 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 430
#2;

verify(ir === 'b1111, "Assert 1716 : < ir !== 'b1111 >");	// Vector No: 429
verify(op === 'b11111111, "Assert 1717 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1718 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1719 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 431
#2;

verify(ir === 'b1111, "Assert 1720 : < ir !== 'b1111 >");	// Vector No: 430
verify(op === 'b11111000, "Assert 1721 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1722 : < extop !== 0 >");
verify(addr === 'b00000111111101111111, "Assert 1723 : < addr !== 'b00000111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 432
#2;

verify(ir === 'b1111, "Assert 1724 : < ir !== 'b1111 >");	// Vector No: 431
verify(op === 'b11111000, "Assert 1725 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1726 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1727 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111111111111111111111111111111111:0:0:1111:11111111:0:11111110111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 433
#2;

verify(ir === 'b1111, "Assert 1728 : < ir !== 'b1111 >");	// Vector No: 432
verify(op === 'b11111111, "Assert 1729 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1730 : < extop !== 0 >");
verify(addr === 'b11111110111111111111, "Assert 1731 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 434
#2;

verify(ir === 'b1111, "Assert 1732 : < ir !== 'b1111 >");	// Vector No: 433
verify(op === 'b11111111, "Assert 1733 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1734 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1735 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 435
#2;

verify(ir === 'b1111, "Assert 1736 : < ir !== 'b1111 >");	// Vector No: 434
verify(op === 'b11111000, "Assert 1737 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1738 : < extop !== 0 >");
verify(addr === 'b00000111111011111111, "Assert 1739 : < addr !== 'b00000111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 436
#2;

verify(ir === 'b1111, "Assert 1740 : < ir !== 'b1111 >");	// Vector No: 435
verify(op === 'b11111000, "Assert 1741 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1742 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1743 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111111111111111111111111111111111:0:0:1111:11111111:0:11111101111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 437
#2;

verify(ir === 'b1111, "Assert 1744 : < ir !== 'b1111 >");	// Vector No: 436
verify(op === 'b11111111, "Assert 1745 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1746 : < extop !== 0 >");
verify(addr === 'b11111101111111111111, "Assert 1747 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 438
#2;

verify(ir === 'b1111, "Assert 1748 : < ir !== 'b1111 >");	// Vector No: 437
verify(op === 'b11111111, "Assert 1749 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1750 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1751 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111110111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 439
#2;

verify(ir === 'b1111, "Assert 1752 : < ir !== 'b1111 >");	// Vector No: 438
verify(op === 'b11111000, "Assert 1753 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1754 : < extop !== 0 >");
verify(addr === 'b00000111110111111111, "Assert 1755 : < addr !== 'b00000111110111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 440
#2;

verify(ir === 'b1111, "Assert 1756 : < ir !== 'b1111 >");	// Vector No: 439
verify(op === 'b11111000, "Assert 1757 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1758 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1759 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111111111111111111111111111111111:0:0:1111:11111111:0:11111011111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 441
#2;

verify(ir === 'b1111, "Assert 1760 : < ir !== 'b1111 >");	// Vector No: 440
verify(op === 'b11111111, "Assert 1761 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1762 : < extop !== 0 >");
verify(addr === 'b11111011111111111111, "Assert 1763 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 442
#2;

verify(ir === 'b1111, "Assert 1764 : < ir !== 'b1111 >");	// Vector No: 441
verify(op === 'b11111111, "Assert 1765 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1766 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1767 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111101111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 443
#2;

verify(ir === 'b1111, "Assert 1768 : < ir !== 'b1111 >");	// Vector No: 442
verify(op === 'b11111000, "Assert 1769 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1770 : < extop !== 0 >");
verify(addr === 'b00000111101111111111, "Assert 1771 : < addr !== 'b00000111101111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 444
#2;

verify(ir === 'b1111, "Assert 1772 : < ir !== 'b1111 >");	// Vector No: 443
verify(op === 'b11111000, "Assert 1773 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1774 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1775 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111111111111111111111111111111111:0:0:1111:11111111:0:11110111111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 445
#2;

verify(ir === 'b1111, "Assert 1776 : < ir !== 'b1111 >");	// Vector No: 444
verify(op === 'b11111111, "Assert 1777 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1778 : < extop !== 0 >");
verify(addr === 'b11110111111111111111, "Assert 1779 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 446
#2;

verify(ir === 'b1111, "Assert 1780 : < ir !== 'b1111 >");	// Vector No: 445
verify(op === 'b11111111, "Assert 1781 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1782 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1783 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111011111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 447
#2;

verify(ir === 'b1111, "Assert 1784 : < ir !== 'b1111 >");	// Vector No: 446
verify(op === 'b11111000, "Assert 1785 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1786 : < extop !== 0 >");
verify(addr === 'b00000111011111111111, "Assert 1787 : < addr !== 'b00000111011111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 448
#2;

verify(ir === 'b1111, "Assert 1788 : < ir !== 'b1111 >");	// Vector No: 447
verify(op === 'b11111000, "Assert 1789 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1790 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1791 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111111111111111111111111111111111:0:0:1111:11111111:0:11101111111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 449
#2;

verify(ir === 'b1111, "Assert 1792 : < ir !== 'b1111 >");	// Vector No: 448
verify(op === 'b11111111, "Assert 1793 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1794 : < extop !== 0 >");
verify(addr === 'b11101111111111111111, "Assert 1795 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 450
#2;

verify(ir === 'b1111, "Assert 1796 : < ir !== 'b1111 >");	// Vector No: 449
verify(op === 'b11111111, "Assert 1797 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1798 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1799 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000110111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 451
#2;

verify(ir === 'b1111, "Assert 1800 : < ir !== 'b1111 >");	// Vector No: 450
verify(op === 'b11111000, "Assert 1801 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1802 : < extop !== 0 >");
verify(addr === 'b00000110111111111111, "Assert 1803 : < addr !== 'b00000110111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 452
#2;

verify(ir === 'b1111, "Assert 1804 : < ir !== 'b1111 >");	// Vector No: 451
verify(op === 'b11111000, "Assert 1805 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1806 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1807 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111111111111111111111111111111111:0:0:1111:11111111:0:11011111111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 453
#2;

verify(ir === 'b1111, "Assert 1808 : < ir !== 'b1111 >");	// Vector No: 452
verify(op === 'b11111111, "Assert 1809 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1810 : < extop !== 0 >");
verify(addr === 'b11011111111111111111, "Assert 1811 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 454
#2;

verify(ir === 'b1111, "Assert 1812 : < ir !== 'b1111 >");	// Vector No: 453
verify(op === 'b11111111, "Assert 1813 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1814 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1815 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000101111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 455
#2;

verify(ir === 'b1111, "Assert 1816 : < ir !== 'b1111 >");	// Vector No: 454
verify(op === 'b11111000, "Assert 1817 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1818 : < extop !== 0 >");
verify(addr === 'b00000101111111111111, "Assert 1819 : < addr !== 'b00000101111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 456
#2;

verify(ir === 'b1111, "Assert 1820 : < ir !== 'b1111 >");	// Vector No: 455
verify(op === 'b11111000, "Assert 1821 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1822 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1823 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111111111111111111111111111111111:0:0:1111:11111111:0:10111111111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 457
#2;

verify(ir === 'b1111, "Assert 1824 : < ir !== 'b1111 >");	// Vector No: 456
verify(op === 'b11111111, "Assert 1825 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1826 : < extop !== 0 >");
verify(addr === 'b10111111111111111111, "Assert 1827 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 458
#2;

verify(ir === 'b1111, "Assert 1828 : < ir !== 'b1111 >");	// Vector No: 457
verify(op === 'b11111111, "Assert 1829 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1830 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1831 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 459
#2;

verify(ir === 'b1111, "Assert 1832 : < ir !== 'b1111 >");	// Vector No: 458
verify(op === 'b11111000, "Assert 1833 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1834 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 1835 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 460
#2;

verify(ir === 'b1111, "Assert 1836 : < ir !== 'b1111 >");	// Vector No: 459
verify(op === 'b11111000, "Assert 1837 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1838 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1839 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111111111111111111111111111111111:0:0:1111:11111111:0:01111111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 461
#2;

verify(ir === 'b1111, "Assert 1840 : < ir !== 'b1111 >");	// Vector No: 460
verify(op === 'b11111111, "Assert 1841 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1842 : < extop !== 0 >");
verify(addr === 'b01111111111111111111, "Assert 1843 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 462
#2;

verify(ir === 'b1111, "Assert 1844 : < ir !== 'b1111 >");	// Vector No: 461
verify(op === 'b11111111, "Assert 1845 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1846 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1847 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111111111111111111111111111111111:1:0:1111:11110000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 463
#2;

verify(ir === 'b1111, "Assert 1848 : < ir !== 'b1111 >");	// Vector No: 462
verify(op === 'b11110000, "Assert 1849 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 1850 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1851 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 464
#2;

verify(ir === 'b1111, "Assert 1852 : < ir !== 'b1111 >");	// Vector No: 463
verify(op === 'b11111000, "Assert 1853 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1854 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1855 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111111111111111111111111111111111:0:0:1111:11111110:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 465
#2;

verify(ir === 'b1111, "Assert 1856 : < ir !== 'b1111 >");	// Vector No: 464
verify(op === 'b11111110, "Assert 1857 : < op !== 'b11111110 >");
verify(extop === 0, "Assert 1858 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1859 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 466
#2;

verify(ir === 'b1111, "Assert 1860 : < ir !== 'b1111 >");	// Vector No: 465
verify(op === 'b11111111, "Assert 1861 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1862 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1863 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111111111111111111111111111111111:1:0:1111:11101000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 467
#2;

verify(ir === 'b1111, "Assert 1864 : < ir !== 'b1111 >");	// Vector No: 466
verify(op === 'b11101000, "Assert 1865 : < op !== 'b11101000 >");
verify(extop === 0, "Assert 1866 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1867 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 468
#2;

verify(ir === 'b1111, "Assert 1868 : < ir !== 'b1111 >");	// Vector No: 467
verify(op === 'b11111000, "Assert 1869 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1870 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1871 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111111111111111111111111111111111:0:0:1111:11111101:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 469
#2;

verify(ir === 'b1111, "Assert 1872 : < ir !== 'b1111 >");	// Vector No: 468
verify(op === 'b11111101, "Assert 1873 : < op !== 'b11111101 >");
verify(extop === 0, "Assert 1874 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1875 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 470
#2;

verify(ir === 'b1111, "Assert 1876 : < ir !== 'b1111 >");	// Vector No: 469
verify(op === 'b11111111, "Assert 1877 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1878 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1879 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111111111111111111111111111111111:1:0:1111:11011000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 471
#2;

verify(ir === 'b1111, "Assert 1880 : < ir !== 'b1111 >");	// Vector No: 470
verify(op === 'b11011000, "Assert 1881 : < op !== 'b11011000 >");
verify(extop === 0, "Assert 1882 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1883 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 472
#2;

verify(ir === 'b1111, "Assert 1884 : < ir !== 'b1111 >");	// Vector No: 471
verify(op === 'b11111000, "Assert 1885 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1886 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1887 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111111111111111111111111111111111:0:0:1111:11111011:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 473
#2;

verify(ir === 'b1111, "Assert 1888 : < ir !== 'b1111 >");	// Vector No: 472
verify(op === 'b11111011, "Assert 1889 : < op !== 'b11111011 >");
verify(extop === 0, "Assert 1890 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1891 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 474
#2;

verify(ir === 'b1111, "Assert 1892 : < ir !== 'b1111 >");	// Vector No: 473
verify(op === 'b11111111, "Assert 1893 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1894 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1895 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111111111111111111111111111111111:1:0:1111:10111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 475
#2;

verify(ir === 'b1111, "Assert 1896 : < ir !== 'b1111 >");	// Vector No: 474
verify(op === 'b10111000, "Assert 1897 : < op !== 'b10111000 >");
verify(extop === 0, "Assert 1898 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1899 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 476
#2;

verify(ir === 'b1111, "Assert 1900 : < ir !== 'b1111 >");	// Vector No: 475
verify(op === 'b11111000, "Assert 1901 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1902 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1903 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111111111111111111111111111111111:0:0:1111:11110111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 477
#2;

verify(ir === 'b1111, "Assert 1904 : < ir !== 'b1111 >");	// Vector No: 476
verify(op === 'b11110111, "Assert 1905 : < op !== 'b11110111 >");
verify(extop === 0, "Assert 1906 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1907 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 478
#2;

verify(ir === 'b1111, "Assert 1908 : < ir !== 'b1111 >");	// Vector No: 477
verify(op === 'b11111111, "Assert 1909 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1910 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1911 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111111111111111111111111111111111:1:0:1111:01111111:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 479
#2;

verify(ir === 'b1111, "Assert 1912 : < ir !== 'b1111 >");	// Vector No: 478
verify(op === 'b01111111, "Assert 1913 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 1914 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1915 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 480
#2;

verify(ir === 'b1111, "Assert 1916 : < ir !== 'b1111 >");	// Vector No: 479
verify(op === 'b11111000, "Assert 1917 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1918 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1919 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111111111111111111111111111111111:0:0:1111:11101111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 481
#2;

verify(ir === 'b1111, "Assert 1920 : < ir !== 'b1111 >");	// Vector No: 480
verify(op === 'b11101111, "Assert 1921 : < op !== 'b11101111 >");
verify(extop === 0, "Assert 1922 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1923 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 482
#2;

verify(ir === 'b1111, "Assert 1924 : < ir !== 'b1111 >");	// Vector No: 481
verify(op === 'b11111111, "Assert 1925 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1926 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1927 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111111111111111111111111111111111:1:0:1110:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 483
#2;

verify(ir === 'b1110, "Assert 1928 : < ir !== 'b1110 >");	// Vector No: 482
verify(op === 'b11111000, "Assert 1929 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1930 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1931 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 484
#2;

verify(ir === 'b1111, "Assert 1932 : < ir !== 'b1111 >");	// Vector No: 483
verify(op === 'b11111000, "Assert 1933 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1934 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1935 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111111111111111111111111111111111:0:0:1111:11011111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 485
#2;

verify(ir === 'b1111, "Assert 1936 : < ir !== 'b1111 >");	// Vector No: 484
verify(op === 'b11011111, "Assert 1937 : < op !== 'b11011111 >");
verify(extop === 0, "Assert 1938 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1939 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 486
#2;

verify(ir === 'b1111, "Assert 1940 : < ir !== 'b1111 >");	// Vector No: 485
verify(op === 'b11111111, "Assert 1941 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1942 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1943 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111111111111111111111111111111111:1:0:1101:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 487
#2;

verify(ir === 'b1101, "Assert 1944 : < ir !== 'b1101 >");	// Vector No: 486
verify(op === 'b11111000, "Assert 1945 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1946 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1947 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 488
#2;

verify(ir === 'b1111, "Assert 1948 : < ir !== 'b1111 >");	// Vector No: 487
verify(op === 'b11111000, "Assert 1949 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1950 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1951 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111111111111111111111111111111111:0:0:1111:10111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 489
#2;

verify(ir === 'b1111, "Assert 1952 : < ir !== 'b1111 >");	// Vector No: 488
verify(op === 'b10111111, "Assert 1953 : < op !== 'b10111111 >");
verify(extop === 0, "Assert 1954 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1955 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 490
#2;

verify(ir === 'b1111, "Assert 1956 : < ir !== 'b1111 >");	// Vector No: 489
verify(op === 'b11111111, "Assert 1957 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1958 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1959 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 491
#2;

verify(ir === 'b1011, "Assert 1960 : < ir !== 'b1011 >");	// Vector No: 490
verify(op === 'b11111000, "Assert 1961 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1962 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1963 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 492
#2;

verify(ir === 'b1111, "Assert 1964 : < ir !== 'b1111 >");	// Vector No: 491
verify(op === 'b11111000, "Assert 1965 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1966 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1967 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111111111111111111111111111111111:0:0:1111:01111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 493
#2;

verify(ir === 'b1111, "Assert 1968 : < ir !== 'b1111 >");	// Vector No: 492
verify(op === 'b01111111, "Assert 1969 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 1970 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1971 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 494
#2;

verify(ir === 'b1111, "Assert 1972 : < ir !== 'b1111 >");	// Vector No: 493
verify(op === 'b11111111, "Assert 1973 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1974 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1975 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 495
#2;

verify(ir === 'b1111, "Assert 1976 : < ir !== 'b1111 >");	// Vector No: 494
verify(op === 'b11111000, "Assert 1977 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1978 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1979 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 496
#2;

verify(ir === 'b1111, "Assert 1980 : < ir !== 'b1111 >");	// Vector No: 495
verify(op === 'b11111000, "Assert 1981 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1982 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1983 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111111111111111111111111111111111:0:0:1110:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 497
#2;

verify(ir === 'b1110, "Assert 1984 : < ir !== 'b1110 >");	// Vector No: 496
verify(op === 'b11111111, "Assert 1985 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1986 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1987 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 498
#2;

verify(ir === 'b1111, "Assert 1988 : < ir !== 'b1111 >");	// Vector No: 497
verify(op === 'b11111111, "Assert 1989 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 1990 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 1991 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 499
#2;

verify(ir === 'b1111, "Assert 1992 : < ir !== 'b1111 >");	// Vector No: 498
verify(op === 'b11111000, "Assert 1993 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1994 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1995 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 500
#2;

verify(ir === 'b1111, "Assert 1996 : < ir !== 'b1111 >");	// Vector No: 499
verify(op === 'b11111000, "Assert 1997 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 1998 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 1999 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111111111111111111111111111111111:0:0:1101:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 501
#2;

verify(ir === 'b1101, "Assert 2000 : < ir !== 'b1101 >");	// Vector No: 500
verify(op === 'b11111111, "Assert 2001 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2002 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2003 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 502
#2;

verify(ir === 'b1111, "Assert 2004 : < ir !== 'b1111 >");	// Vector No: 501
verify(op === 'b11111111, "Assert 2005 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2006 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2007 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 503
#2;

verify(ir === 'b1111, "Assert 2008 : < ir !== 'b1111 >");	// Vector No: 502
verify(op === 'b11111000, "Assert 2009 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2010 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2011 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 504
#2;

verify(ir === 'b1111, "Assert 2012 : < ir !== 'b1111 >");	// Vector No: 503
verify(op === 'b11111000, "Assert 2013 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2014 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2015 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111111111111111111111111111111111:0:0:1011:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 505
#2;

verify(ir === 'b1011, "Assert 2016 : < ir !== 'b1011 >");	// Vector No: 504
verify(op === 'b11111111, "Assert 2017 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2018 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2019 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 506
#2;

verify(ir === 'b1111, "Assert 2020 : < ir !== 'b1111 >");	// Vector No: 505
verify(op === 'b11111111, "Assert 2021 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2022 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2023 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111111111111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 507
#2;

verify(ir === 'b1111, "Assert 2024 : < ir !== 'b1111 >");	// Vector No: 506
verify(op === 'b11111000, "Assert 2025 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2026 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2027 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 508
#2;

verify(ir === 'b1111, "Assert 2028 : < ir !== 'b1111 >");	// Vector No: 507
verify(op === 'b11111000, "Assert 2029 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2030 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2031 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111111111111111111111111111111111:0:0:0111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 509
#2;

verify(ir === 'b0111, "Assert 2032 : < ir !== 'b0111 >");	// Vector No: 508
verify(op === 'b11111111, "Assert 2033 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2034 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2035 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 510
#2;

verify(ir === 'b1111, "Assert 2036 : < ir !== 'b1111 >");	// Vector No: 509
verify(op === 'b11111111, "Assert 2037 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 2038 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 2039 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111111111111111111111111111111111:1:0:0111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 511
#2;

verify(ir === 'b0111, "Assert 2040 : < ir !== 'b0111 >");	// Vector No: 510
verify(op === 'b11111000, "Assert 2041 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2042 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2043 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 512
#2;

verify(ir === 'b1111, "Assert 2044 : < ir !== 'b1111 >");	// Vector No: 511
verify(op === 'b11111000, "Assert 2045 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 2046 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 2047 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000001:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 513
#2;

verify(ir === 'b0000, "Assert 2048 : < ir !== 'b0000 >");	// Vector No: 512
verify(op === 'b00000000, "Assert 2049 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2050 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2051 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000001:0:1:1000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 514
#2;

verify(ir === 'b1000, "Assert 2052 : < ir !== 'b1000 >");	// Vector No: 513
verify(op === 'b00000000, "Assert 2053 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2054 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 2055 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000001:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 515
#2;

verify(ir === 'b0000, "Assert 2056 : < ir !== 'b0000 >");	// Vector No: 514
verify(op === 'b00000000, "Assert 2057 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2058 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2059 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000001:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 516
#2;

verify(ir === 'b0000, "Assert 2060 : < ir !== 'b0000 >");	// Vector No: 515
verify(op === 'b00000000, "Assert 2061 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2062 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2063 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000010:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 517
#2;

verify(ir === 'b0000, "Assert 2064 : < ir !== 'b0000 >");	// Vector No: 516
verify(op === 'b00000000, "Assert 2065 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2066 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2067 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000010:0:1:1000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 518
#2;

verify(ir === 'b1000, "Assert 2068 : < ir !== 'b1000 >");	// Vector No: 517
verify(op === 'b00000000, "Assert 2069 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2070 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 2071 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000010:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 519
#2;

verify(ir === 'b0000, "Assert 2072 : < ir !== 'b0000 >");	// Vector No: 518
verify(op === 'b00000000, "Assert 2073 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2074 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2075 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000010:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 520
#2;

verify(ir === 'b0000, "Assert 2076 : < ir !== 'b0000 >");	// Vector No: 519
verify(op === 'b00000000, "Assert 2077 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2078 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2079 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000100:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 521
#2;

verify(ir === 'b0000, "Assert 2080 : < ir !== 'b0000 >");	// Vector No: 520
verify(op === 'b00000000, "Assert 2081 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2082 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2083 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000100:0:1:1000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 522
#2;

verify(ir === 'b1000, "Assert 2084 : < ir !== 'b1000 >");	// Vector No: 521
verify(op === 'b00000000, "Assert 2085 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2086 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 2087 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000100:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 523
#2;

verify(ir === 'b0000, "Assert 2088 : < ir !== 'b0000 >");	// Vector No: 522
verify(op === 'b00000000, "Assert 2089 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2090 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2091 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000000100:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 524
#2;

verify(ir === 'b0000, "Assert 2092 : < ir !== 'b0000 >");	// Vector No: 523
verify(op === 'b00000000, "Assert 2093 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2094 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2095 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000001000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 525
#2;

verify(ir === 'b0000, "Assert 2096 : < ir !== 'b0000 >");	// Vector No: 524
verify(op === 'b00000000, "Assert 2097 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2098 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2099 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000001000:0:1:1000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 526
#2;

verify(ir === 'b1000, "Assert 2100 : < ir !== 'b1000 >");	// Vector No: 525
verify(op === 'b00000000, "Assert 2101 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2102 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 2103 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000001000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 527
#2;

verify(ir === 'b0000, "Assert 2104 : < ir !== 'b0000 >");	// Vector No: 526
verify(op === 'b00000000, "Assert 2105 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2106 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2107 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000001000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 528
#2;

verify(ir === 'b0000, "Assert 2108 : < ir !== 'b0000 >");	// Vector No: 527
verify(op === 'b00000000, "Assert 2109 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2110 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2111 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000010000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 529
#2;

verify(ir === 'b0000, "Assert 2112 : < ir !== 'b0000 >");	// Vector No: 528
verify(op === 'b00000000, "Assert 2113 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2114 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2115 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000010000:0:1:1000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 530
#2;

verify(ir === 'b1000, "Assert 2116 : < ir !== 'b1000 >");	// Vector No: 529
verify(op === 'b00000000, "Assert 2117 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2118 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 2119 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000010000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 531
#2;

verify(ir === 'b0000, "Assert 2120 : < ir !== 'b0000 >");	// Vector No: 530
verify(op === 'b00000000, "Assert 2121 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2122 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2123 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000010000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 532
#2;

verify(ir === 'b0000, "Assert 2124 : < ir !== 'b0000 >");	// Vector No: 531
verify(op === 'b00000000, "Assert 2125 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2126 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2127 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000100000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 533
#2;

verify(ir === 'b0000, "Assert 2128 : < ir !== 'b0000 >");	// Vector No: 532
verify(op === 'b00000000, "Assert 2129 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2130 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2131 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000100000:0:1:1000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 534
#2;

verify(ir === 'b1000, "Assert 2132 : < ir !== 'b1000 >");	// Vector No: 533
verify(op === 'b00000000, "Assert 2133 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2134 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 2135 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000100000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 535
#2;

verify(ir === 'b0000, "Assert 2136 : < ir !== 'b0000 >");	// Vector No: 534
verify(op === 'b00000000, "Assert 2137 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2138 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2139 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000000100000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 536
#2;

verify(ir === 'b0000, "Assert 2140 : < ir !== 'b0000 >");	// Vector No: 535
verify(op === 'b00000000, "Assert 2141 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2142 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2143 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000001000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 537
#2;

verify(ir === 'b0000, "Assert 2144 : < ir !== 'b0000 >");	// Vector No: 536
verify(op === 'b00000000, "Assert 2145 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2146 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2147 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000001000000:0:1:1000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 538
#2;

verify(ir === 'b1000, "Assert 2148 : < ir !== 'b1000 >");	// Vector No: 537
verify(op === 'b00000000, "Assert 2149 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2150 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 2151 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000001000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 539
#2;

verify(ir === 'b0000, "Assert 2152 : < ir !== 'b0000 >");	// Vector No: 538
verify(op === 'b00000000, "Assert 2153 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2154 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2155 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000001000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 540
#2;

verify(ir === 'b0000, "Assert 2156 : < ir !== 'b0000 >");	// Vector No: 539
verify(op === 'b00000000, "Assert 2157 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2158 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2159 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000010000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 541
#2;

verify(ir === 'b0000, "Assert 2160 : < ir !== 'b0000 >");	// Vector No: 540
verify(op === 'b00000000, "Assert 2161 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2162 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2163 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000010000000:0:1:1000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 542
#2;

verify(ir === 'b1000, "Assert 2164 : < ir !== 'b1000 >");	// Vector No: 541
verify(op === 'b00000000, "Assert 2165 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2166 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 2167 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000010000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 543
#2;

verify(ir === 'b0000, "Assert 2168 : < ir !== 'b0000 >");	// Vector No: 542
verify(op === 'b00000000, "Assert 2169 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2170 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2171 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000010000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 544
#2;

verify(ir === 'b0000, "Assert 2172 : < ir !== 'b0000 >");	// Vector No: 543
verify(op === 'b00000000, "Assert 2173 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2174 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2175 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000100000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 545
#2;

verify(ir === 'b0000, "Assert 2176 : < ir !== 'b0000 >");	// Vector No: 544
verify(op === 'b00000000, "Assert 2177 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2178 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2179 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000100000000:0:1:1000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 546
#2;

verify(ir === 'b1000, "Assert 2180 : < ir !== 'b1000 >");	// Vector No: 545
verify(op === 'b00000000, "Assert 2181 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2182 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 2183 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000100000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 547
#2;

verify(ir === 'b0000, "Assert 2184 : < ir !== 'b0000 >");	// Vector No: 546
verify(op === 'b00000000, "Assert 2185 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2186 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2187 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000000100000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 548
#2;

verify(ir === 'b0000, "Assert 2188 : < ir !== 'b0000 >");	// Vector No: 547
verify(op === 'b00000000, "Assert 2189 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2190 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2191 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000001000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 549
#2;

verify(ir === 'b0000, "Assert 2192 : < ir !== 'b0000 >");	// Vector No: 548
verify(op === 'b00000000, "Assert 2193 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2194 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2195 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000001000000000:0:1:1000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 550
#2;

verify(ir === 'b1000, "Assert 2196 : < ir !== 'b1000 >");	// Vector No: 549
verify(op === 'b00000000, "Assert 2197 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2198 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 2199 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000001000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 551
#2;

verify(ir === 'b0000, "Assert 2200 : < ir !== 'b0000 >");	// Vector No: 550
verify(op === 'b00000000, "Assert 2201 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2202 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2203 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000001000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 552
#2;

verify(ir === 'b0000, "Assert 2204 : < ir !== 'b0000 >");	// Vector No: 551
verify(op === 'b00000000, "Assert 2205 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2206 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2207 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000010000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 553
#2;

verify(ir === 'b0000, "Assert 2208 : < ir !== 'b0000 >");	// Vector No: 552
verify(op === 'b00000000, "Assert 2209 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2210 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2211 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000010000000000:0:1:1000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 554
#2;

verify(ir === 'b1000, "Assert 2212 : < ir !== 'b1000 >");	// Vector No: 553
verify(op === 'b00000000, "Assert 2213 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2214 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 2215 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000010000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 555
#2;

verify(ir === 'b0000, "Assert 2216 : < ir !== 'b0000 >");	// Vector No: 554
verify(op === 'b00000000, "Assert 2217 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2218 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2219 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000010000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 556
#2;

verify(ir === 'b0000, "Assert 2220 : < ir !== 'b0000 >");	// Vector No: 555
verify(op === 'b00000000, "Assert 2221 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2222 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2223 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000100000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 557
#2;

verify(ir === 'b0000, "Assert 2224 : < ir !== 'b0000 >");	// Vector No: 556
verify(op === 'b00000000, "Assert 2225 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2226 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2227 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000100000000000:0:1:1000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 558
#2;

verify(ir === 'b1000, "Assert 2228 : < ir !== 'b1000 >");	// Vector No: 557
verify(op === 'b00000000, "Assert 2229 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2230 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 2231 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000100000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 559
#2;

verify(ir === 'b0000, "Assert 2232 : < ir !== 'b0000 >");	// Vector No: 558
verify(op === 'b00000000, "Assert 2233 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2234 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2235 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000000100000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 560
#2;

verify(ir === 'b0000, "Assert 2236 : < ir !== 'b0000 >");	// Vector No: 559
verify(op === 'b00000000, "Assert 2237 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2238 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2239 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000001000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 561
#2;

verify(ir === 'b0000, "Assert 2240 : < ir !== 'b0000 >");	// Vector No: 560
verify(op === 'b00000000, "Assert 2241 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2242 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2243 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000001000000000000:0:1:1000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 562
#2;

verify(ir === 'b1000, "Assert 2244 : < ir !== 'b1000 >");	// Vector No: 561
verify(op === 'b00000000, "Assert 2245 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2246 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 2247 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000001000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 563
#2;

verify(ir === 'b0000, "Assert 2248 : < ir !== 'b0000 >");	// Vector No: 562
verify(op === 'b00000000, "Assert 2249 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2250 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2251 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000001000000000000:1:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 564
#2;

verify(ir === 'b0000, "Assert 2252 : < ir !== 'b0000 >");	// Vector No: 563
verify(op === 'b00000000, "Assert 2253 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2254 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 2255 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000010000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 565
#2;

verify(ir === 'b0000, "Assert 2256 : < ir !== 'b0000 >");	// Vector No: 564
verify(op === 'b00000000, "Assert 2257 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2258 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2259 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000010000000000000:0:1:1000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 566
#2;

verify(ir === 'b1000, "Assert 2260 : < ir !== 'b1000 >");	// Vector No: 565
verify(op === 'b00000000, "Assert 2261 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2262 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 2263 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000010000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 567
#2;

verify(ir === 'b0000, "Assert 2264 : < ir !== 'b0000 >");	// Vector No: 566
verify(op === 'b00000000, "Assert 2265 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2266 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2267 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000010000000000000:1:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 568
#2;

verify(ir === 'b0000, "Assert 2268 : < ir !== 'b0000 >");	// Vector No: 567
verify(op === 'b00000000, "Assert 2269 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2270 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 2271 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000100000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 569
#2;

verify(ir === 'b0000, "Assert 2272 : < ir !== 'b0000 >");	// Vector No: 568
verify(op === 'b00000000, "Assert 2273 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2274 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2275 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000100000000000000:0:1:1000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 570
#2;

verify(ir === 'b1000, "Assert 2276 : < ir !== 'b1000 >");	// Vector No: 569
verify(op === 'b00000000, "Assert 2277 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2278 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 2279 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000100000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 571
#2;

verify(ir === 'b0000, "Assert 2280 : < ir !== 'b0000 >");	// Vector No: 570
verify(op === 'b00000000, "Assert 2281 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2282 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2283 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000000100000000000000:1:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000000100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 572
#2;

verify(ir === 'b0000, "Assert 2284 : < ir !== 'b0000 >");	// Vector No: 571
verify(op === 'b00000000, "Assert 2285 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2286 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 2287 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000001000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000001000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 573
#2;

verify(ir === 'b0000, "Assert 2288 : < ir !== 'b0000 >");	// Vector No: 572
verify(op === 'b00000000, "Assert 2289 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2290 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2291 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000001000000000000000:0:1:1000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000001000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 574
#2;

verify(ir === 'b1000, "Assert 2292 : < ir !== 'b1000 >");	// Vector No: 573
verify(op === 'b00000000, "Assert 2293 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2294 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 2295 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000001000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000001000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 575
#2;

verify(ir === 'b0000, "Assert 2296 : < ir !== 'b0000 >");	// Vector No: 574
verify(op === 'b00000000, "Assert 2297 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2298 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2299 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000001000000000000000:1:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000001000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 576
#2;

verify(ir === 'b0000, "Assert 2300 : < ir !== 'b0000 >");	// Vector No: 575
verify(op === 'b00000000, "Assert 2301 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2302 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 2303 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000010000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000010000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 577
#2;

verify(ir === 'b0000, "Assert 2304 : < ir !== 'b0000 >");	// Vector No: 576
verify(op === 'b00000000, "Assert 2305 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2306 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2307 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000010000000000000000:0:1:1000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000010000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 578
#2;

verify(ir === 'b1000, "Assert 2308 : < ir !== 'b1000 >");	// Vector No: 577
verify(op === 'b00000000, "Assert 2309 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2310 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 2311 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000010000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000010000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 579
#2;

verify(ir === 'b0000, "Assert 2312 : < ir !== 'b0000 >");	// Vector No: 578
verify(op === 'b00000000, "Assert 2313 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2314 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2315 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000010000000000000000:1:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000010000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 580
#2;

verify(ir === 'b0000, "Assert 2316 : < ir !== 'b0000 >");	// Vector No: 579
verify(op === 'b00000000, "Assert 2317 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2318 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 2319 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000100000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000100000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 581
#2;

verify(ir === 'b0000, "Assert 2320 : < ir !== 'b0000 >");	// Vector No: 580
verify(op === 'b00000000, "Assert 2321 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2322 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2323 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000100000000000000000:0:1:1000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000100000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 582
#2;

verify(ir === 'b1000, "Assert 2324 : < ir !== 'b1000 >");	// Vector No: 581
verify(op === 'b00000000, "Assert 2325 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2326 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 2327 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000100000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000100000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 583
#2;

verify(ir === 'b0000, "Assert 2328 : < ir !== 'b0000 >");	// Vector No: 582
verify(op === 'b00000000, "Assert 2329 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2330 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2331 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000000100000000000000000:1:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000000100000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 584
#2;

verify(ir === 'b0000, "Assert 2332 : < ir !== 'b0000 >");	// Vector No: 583
verify(op === 'b00000000, "Assert 2333 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2334 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 2335 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000001000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000001000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 585
#2;

verify(ir === 'b0000, "Assert 2336 : < ir !== 'b0000 >");	// Vector No: 584
verify(op === 'b00000000, "Assert 2337 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2338 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2339 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000001000000000000000000:0:1:1000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000001000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 586
#2;

verify(ir === 'b1000, "Assert 2340 : < ir !== 'b1000 >");	// Vector No: 585
verify(op === 'b00000000, "Assert 2341 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2342 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 2343 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000001000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000001000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 587
#2;

verify(ir === 'b0000, "Assert 2344 : < ir !== 'b0000 >");	// Vector No: 586
verify(op === 'b00000000, "Assert 2345 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2346 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2347 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000001000000000000000000:1:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000001000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 588
#2;

verify(ir === 'b0000, "Assert 2348 : < ir !== 'b0000 >");	// Vector No: 587
verify(op === 'b00000000, "Assert 2349 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2350 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 2351 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000010000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000010000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 589
#2;

verify(ir === 'b0000, "Assert 2352 : < ir !== 'b0000 >");	// Vector No: 588
verify(op === 'b00000000, "Assert 2353 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2354 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2355 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000010000000000000000000:0:1:1000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000010000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 590
#2;

verify(ir === 'b1000, "Assert 2356 : < ir !== 'b1000 >");	// Vector No: 589
verify(op === 'b00000000, "Assert 2357 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2358 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 2359 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000010000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000010000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 591
#2;

verify(ir === 'b0000, "Assert 2360 : < ir !== 'b0000 >");	// Vector No: 590
verify(op === 'b00000000, "Assert 2361 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2362 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2363 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000010000000000000000000:1:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000010000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 592
#2;

verify(ir === 'b0000, "Assert 2364 : < ir !== 'b0000 >");	// Vector No: 591
verify(op === 'b00000000, "Assert 2365 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2366 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 2367 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 593
#2;

verify(ir === 'b0000, "Assert 2368 : < ir !== 'b0000 >");	// Vector No: 592
verify(op === 'b00000000, "Assert 2369 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2370 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2371 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000100000000000000000000:0:1:1000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 594
#2;

verify(ir === 'b1000, "Assert 2372 : < ir !== 'b1000 >");	// Vector No: 593
verify(op === 'b00000001, "Assert 2373 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 2374 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2375 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 595
#2;

verify(ir === 'b0000, "Assert 2376 : < ir !== 'b0000 >");	// Vector No: 594
verify(op === 'b00000000, "Assert 2377 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2378 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2379 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000000100000000000000000000:1:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000000100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 596
#2;

verify(ir === 'b0000, "Assert 2380 : < ir !== 'b0000 >");	// Vector No: 595
verify(op === 'b00000000, "Assert 2381 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2382 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 2383 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000001000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000001000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 597
#2;

verify(ir === 'b0000, "Assert 2384 : < ir !== 'b0000 >");	// Vector No: 596
verify(op === 'b00000000, "Assert 2385 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2386 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2387 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000001000000000000000000000:0:1:1000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000001000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 598
#2;

verify(ir === 'b1000, "Assert 2388 : < ir !== 'b1000 >");	// Vector No: 597
verify(op === 'b00000010, "Assert 2389 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 2390 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2391 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000001000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000001000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 599
#2;

verify(ir === 'b0000, "Assert 2392 : < ir !== 'b0000 >");	// Vector No: 598
verify(op === 'b00000000, "Assert 2393 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2394 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2395 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000001000000000000000000000:1:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000001000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 600
#2;

verify(ir === 'b0000, "Assert 2396 : < ir !== 'b0000 >");	// Vector No: 599
verify(op === 'b00000000, "Assert 2397 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2398 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 2399 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000010000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000010000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 601
#2;

verify(ir === 'b0000, "Assert 2400 : < ir !== 'b0000 >");	// Vector No: 600
verify(op === 'b00000000, "Assert 2401 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2402 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2403 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000010000000000000000000000:0:1:1000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000010000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 602
#2;

verify(ir === 'b1000, "Assert 2404 : < ir !== 'b1000 >");	// Vector No: 601
verify(op === 'b00000100, "Assert 2405 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 2406 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2407 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000010000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000010000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 603
#2;

verify(ir === 'b0000, "Assert 2408 : < ir !== 'b0000 >");	// Vector No: 602
verify(op === 'b00000000, "Assert 2409 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2410 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2411 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000010000000000000000000000:1:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000010000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 604
#2;

verify(ir === 'b0000, "Assert 2412 : < ir !== 'b0000 >");	// Vector No: 603
verify(op === 'b00000000, "Assert 2413 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2414 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 2415 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000100000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000100000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 605
#2;

verify(ir === 'b0000, "Assert 2416 : < ir !== 'b0000 >");	// Vector No: 604
verify(op === 'b00000000, "Assert 2417 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2418 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2419 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000100000000000000000000000:0:1:1000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000100000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 606
#2;

verify(ir === 'b1000, "Assert 2420 : < ir !== 'b1000 >");	// Vector No: 605
verify(op === 'b00001000, "Assert 2421 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 2422 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2423 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000100000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000100000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 607
#2;

verify(ir === 'b0000, "Assert 2424 : < ir !== 'b0000 >");	// Vector No: 606
verify(op === 'b00000000, "Assert 2425 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2426 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2427 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000000100000000000000000000000:1:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000000100000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 608
#2;

verify(ir === 'b0000, "Assert 2428 : < ir !== 'b0000 >");	// Vector No: 607
verify(op === 'b00000000, "Assert 2429 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2430 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 2431 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000001000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000001000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 609
#2;

verify(ir === 'b0000, "Assert 2432 : < ir !== 'b0000 >");	// Vector No: 608
verify(op === 'b00000000, "Assert 2433 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2434 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2435 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000001000000000000000000000000:0:1:1000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000001000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 610
#2;

verify(ir === 'b1000, "Assert 2436 : < ir !== 'b1000 >");	// Vector No: 609
verify(op === 'b00010000, "Assert 2437 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 2438 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2439 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000001000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000001000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 611
#2;

verify(ir === 'b0000, "Assert 2440 : < ir !== 'b0000 >");	// Vector No: 610
verify(op === 'b00000000, "Assert 2441 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2442 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2443 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000001000000000000000000000000:1:1:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000001000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 612
#2;

verify(ir === 'b0000, "Assert 2444 : < ir !== 'b0000 >");	// Vector No: 611
verify(op === 'b00000000, "Assert 2445 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2446 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 2447 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000010000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000010000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 613
#2;

verify(ir === 'b0000, "Assert 2448 : < ir !== 'b0000 >");	// Vector No: 612
verify(op === 'b00000000, "Assert 2449 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2450 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2451 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000010000000000000000000000000:0:1:1000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000010000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 614
#2;

verify(ir === 'b1000, "Assert 2452 : < ir !== 'b1000 >");	// Vector No: 613
verify(op === 'b00100000, "Assert 2453 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 2454 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2455 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000010000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000010000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 615
#2;

verify(ir === 'b0000, "Assert 2456 : < ir !== 'b0000 >");	// Vector No: 614
verify(op === 'b00000000, "Assert 2457 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2458 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2459 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000010000000000000000000000000:1:1:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000010000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 616
#2;

verify(ir === 'b0000, "Assert 2460 : < ir !== 'b0000 >");	// Vector No: 615
verify(op === 'b00000000, "Assert 2461 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2462 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 2463 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000100000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000100000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 617
#2;

verify(ir === 'b0000, "Assert 2464 : < ir !== 'b0000 >");	// Vector No: 616
verify(op === 'b00000000, "Assert 2465 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2466 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2467 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000100000000000000000000000000:0:1:1000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000100000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 618
#2;

verify(ir === 'b1000, "Assert 2468 : < ir !== 'b1000 >");	// Vector No: 617
verify(op === 'b01000000, "Assert 2469 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 2470 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2471 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000100000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000100000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 619
#2;

verify(ir === 'b0000, "Assert 2472 : < ir !== 'b0000 >");	// Vector No: 618
verify(op === 'b00000000, "Assert 2473 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2474 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2475 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000100000000000000000000000000:1:1:0000:00001000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000100000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 620
#2;

verify(ir === 'b0000, "Assert 2476 : < ir !== 'b0000 >");	// Vector No: 619
verify(op === 'b00001000, "Assert 2477 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 2478 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 2479 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010001000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010001000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 621
#2;

verify(ir === 'b0000, "Assert 2480 : < ir !== 'b0000 >");	// Vector No: 620
verify(op === 'b00000000, "Assert 2481 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2482 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2483 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010001000000000000000000000000000:0:1:1000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010001000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 622
#2;

verify(ir === 'b1000, "Assert 2484 : < ir !== 'b1000 >");	// Vector No: 621
verify(op === 'b10000000, "Assert 2485 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 2486 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2487 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010001000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010001000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 623
#2;

verify(ir === 'b0000, "Assert 2488 : < ir !== 'b0000 >");	// Vector No: 622
verify(op === 'b00000000, "Assert 2489 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2490 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2491 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010001000000000000000000000000000:1:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010001000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 624
#2;

verify(ir === 'b0000, "Assert 2492 : < ir !== 'b0000 >");	// Vector No: 623
verify(op === 'b00010000, "Assert 2493 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 2494 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2495 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010010000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010010000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 625
#2;

verify(ir === 'b0000, "Assert 2496 : < ir !== 'b0000 >");	// Vector No: 624
verify(op === 'b00000000, "Assert 2497 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2498 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2499 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010010000000000000000000000000000:0:1:1001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010010000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 626
#2;

verify(ir === 'b1001, "Assert 2500 : < ir !== 'b1001 >");	// Vector No: 625
verify(op === 'b00000000, "Assert 2501 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2502 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2503 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010010000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010010000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 627
#2;

verify(ir === 'b0000, "Assert 2504 : < ir !== 'b0000 >");	// Vector No: 626
verify(op === 'b00000000, "Assert 2505 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2506 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2507 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010010000000000000000000000000000:1:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010010000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 628
#2;

verify(ir === 'b0000, "Assert 2508 : < ir !== 'b0000 >");	// Vector No: 627
verify(op === 'b00100000, "Assert 2509 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 2510 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2511 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010100000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010100000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 629
#2;

verify(ir === 'b0000, "Assert 2512 : < ir !== 'b0000 >");	// Vector No: 628
verify(op === 'b00000000, "Assert 2513 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2514 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2515 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010100000000000000000000000000000:0:1:1010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010100000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 630
#2;

verify(ir === 'b1010, "Assert 2516 : < ir !== 'b1010 >");	// Vector No: 629
verify(op === 'b00000000, "Assert 2517 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2518 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2519 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010100000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010100000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 631
#2;

verify(ir === 'b0000, "Assert 2520 : < ir !== 'b0000 >");	// Vector No: 630
verify(op === 'b00000000, "Assert 2521 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2522 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2523 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010100000000000000000000000000000:1:1:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010100000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 632
#2;

verify(ir === 'b0000, "Assert 2524 : < ir !== 'b0000 >");	// Vector No: 631
verify(op === 'b01000000, "Assert 2525 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 2526 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2527 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000011000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000011000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 633
#2;

verify(ir === 'b0000, "Assert 2528 : < ir !== 'b0000 >");	// Vector No: 632
verify(op === 'b00000000, "Assert 2529 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2530 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2531 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000011000000000000000000000000000000:0:1:1100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000011000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 634
#2;

verify(ir === 'b1100, "Assert 2532 : < ir !== 'b1100 >");	// Vector No: 633
verify(op === 'b00000000, "Assert 2533 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2534 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2535 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000011000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000011000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 635
#2;

verify(ir === 'b0000, "Assert 2536 : < ir !== 'b0000 >");	// Vector No: 634
verify(op === 'b00000000, "Assert 2537 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2538 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2539 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000011000000000000000000000000000000:1:1:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000011000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 636
#2;

verify(ir === 'b0000, "Assert 2540 : < ir !== 'b0000 >");	// Vector No: 635
verify(op === 'b10000000, "Assert 2541 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 2542 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2543 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000110000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000110000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 637
#2;

verify(ir === 'b0000, "Assert 2544 : < ir !== 'b0000 >");	// Vector No: 636
verify(op === 'b00000000, "Assert 2545 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2546 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 2547 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000110000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000110000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 638
#2;

verify(ir === 'b1000, "Assert 2548 : < ir !== 'b1000 >");	// Vector No: 637
verify(op === 'b00000000, "Assert 2549 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2550 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2551 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000110000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000110000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 639
#2;

verify(ir === 'b0000, "Assert 2552 : < ir !== 'b0000 >");	// Vector No: 638
verify(op === 'b00000000, "Assert 2553 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2554 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2555 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000110000000000000000000000000000000:1:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000110000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 640
#2;

verify(ir === 'b0001, "Assert 2556 : < ir !== 'b0001 >");	// Vector No: 639
verify(op === 'b00000000, "Assert 2557 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2558 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2559 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000001010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 641
#2;

verify(ir === 'b0000, "Assert 2560 : < ir !== 'b0000 >");	// Vector No: 640
verify(op === 'b00000000, "Assert 2561 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2562 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 2563 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000001010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 642
#2;

verify(ir === 'b1000, "Assert 2564 : < ir !== 'b1000 >");	// Vector No: 641
verify(op === 'b00000000, "Assert 2565 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2566 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2567 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 643
#2;

verify(ir === 'b0000, "Assert 2568 : < ir !== 'b0000 >");	// Vector No: 642
verify(op === 'b00000000, "Assert 2569 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2570 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2571 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001010000000000000000000000000000000:1:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 644
#2;

verify(ir === 'b0010, "Assert 2572 : < ir !== 'b0010 >");	// Vector No: 643
verify(op === 'b00000000, "Assert 2573 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2574 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2575 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000010010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 645
#2;

verify(ir === 'b0000, "Assert 2576 : < ir !== 'b0000 >");	// Vector No: 644
verify(op === 'b00000000, "Assert 2577 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2578 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 2579 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000010010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 646
#2;

verify(ir === 'b1000, "Assert 2580 : < ir !== 'b1000 >");	// Vector No: 645
verify(op === 'b00000000, "Assert 2581 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2582 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2583 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 647
#2;

verify(ir === 'b0000, "Assert 2584 : < ir !== 'b0000 >");	// Vector No: 646
verify(op === 'b00000000, "Assert 2585 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2586 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2587 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010010000000000000000000000000000000:1:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 648
#2;

verify(ir === 'b0100, "Assert 2588 : < ir !== 'b0100 >");	// Vector No: 647
verify(op === 'b00000000, "Assert 2589 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2590 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2591 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 649
#2;

verify(ir === 'b0000, "Assert 2592 : < ir !== 'b0000 >");	// Vector No: 648
verify(op === 'b00000000, "Assert 2593 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2594 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 2595 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 650
#2;

verify(ir === 'b1000, "Assert 2596 : < ir !== 'b1000 >");	// Vector No: 649
verify(op === 'b00000000, "Assert 2597 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2598 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2599 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 651
#2;

verify(ir === 'b0000, "Assert 2600 : < ir !== 'b0000 >");	// Vector No: 650
verify(op === 'b00000000, "Assert 2601 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2602 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2603 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100010000000000000000000000000000000:1:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 652
#2;

verify(ir === 'b1000, "Assert 2604 : < ir !== 'b1000 >");	// Vector No: 651
verify(op === 'b00000000, "Assert 2605 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2606 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2607 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 653
#2;

verify(ir === 'b0000, "Assert 2608 : < ir !== 'b0000 >");	// Vector No: 652
verify(op === 'b00000000, "Assert 2609 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2610 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 2611 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 654
#2;

verify(ir === 'b1000, "Assert 2612 : < ir !== 'b1000 >");	// Vector No: 653
verify(op === 'b00000000, "Assert 2613 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2614 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2615 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000001000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 655
#2;

verify(ir === 'b0000, "Assert 2616 : < ir !== 'b0000 >");	// Vector No: 654
verify(op === 'b00000000, "Assert 2617 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2618 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 2619 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000001000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 656
#2;

verify(ir === 'b0000, "Assert 2620 : < ir !== 'b0000 >");	// Vector No: 655
verify(op === 'b00000000, "Assert 2621 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2622 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2623 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 657
#2;

verify(ir === 'b0000, "Assert 2624 : < ir !== 'b0000 >");	// Vector No: 656
verify(op === 'b00000000, "Assert 2625 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2626 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 2627 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 658
#2;

verify(ir === 'b1000, "Assert 2628 : < ir !== 'b1000 >");	// Vector No: 657
verify(op === 'b00000000, "Assert 2629 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2630 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2631 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000010000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 659
#2;

verify(ir === 'b0000, "Assert 2632 : < ir !== 'b0000 >");	// Vector No: 658
verify(op === 'b00000000, "Assert 2633 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2634 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 2635 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000010000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 660
#2;

verify(ir === 'b0000, "Assert 2636 : < ir !== 'b0000 >");	// Vector No: 659
verify(op === 'b00000000, "Assert 2637 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2638 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2639 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 661
#2;

verify(ir === 'b0000, "Assert 2640 : < ir !== 'b0000 >");	// Vector No: 660
verify(op === 'b00000000, "Assert 2641 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2642 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 2643 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 662
#2;

verify(ir === 'b1000, "Assert 2644 : < ir !== 'b1000 >");	// Vector No: 661
verify(op === 'b00000000, "Assert 2645 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2646 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2647 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000100000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 663
#2;

verify(ir === 'b0000, "Assert 2648 : < ir !== 'b0000 >");	// Vector No: 662
verify(op === 'b00000000, "Assert 2649 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2650 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 2651 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000100000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 664
#2;

verify(ir === 'b0000, "Assert 2652 : < ir !== 'b0000 >");	// Vector No: 663
verify(op === 'b00000000, "Assert 2653 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2654 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2655 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 665
#2;

verify(ir === 'b0000, "Assert 2656 : < ir !== 'b0000 >");	// Vector No: 664
verify(op === 'b00000000, "Assert 2657 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2658 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 2659 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 666
#2;

verify(ir === 'b1000, "Assert 2660 : < ir !== 'b1000 >");	// Vector No: 665
verify(op === 'b00000000, "Assert 2661 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2662 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2663 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 667
#2;

verify(ir === 'b0000, "Assert 2664 : < ir !== 'b0000 >");	// Vector No: 666
verify(op === 'b00000000, "Assert 2665 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2666 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 2667 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 668
#2;

verify(ir === 'b0000, "Assert 2668 : < ir !== 'b0000 >");	// Vector No: 667
verify(op === 'b00000000, "Assert 2669 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2670 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2671 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 669
#2;

verify(ir === 'b0000, "Assert 2672 : < ir !== 'b0000 >");	// Vector No: 668
verify(op === 'b00000000, "Assert 2673 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2674 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 2675 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 670
#2;

verify(ir === 'b1000, "Assert 2676 : < ir !== 'b1000 >");	// Vector No: 669
verify(op === 'b00000000, "Assert 2677 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2678 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2679 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 671
#2;

verify(ir === 'b0000, "Assert 2680 : < ir !== 'b0000 >");	// Vector No: 670
verify(op === 'b00000000, "Assert 2681 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2682 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 2683 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 672
#2;

verify(ir === 'b0000, "Assert 2684 : < ir !== 'b0000 >");	// Vector No: 671
verify(op === 'b00000000, "Assert 2685 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2686 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2687 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 673
#2;

verify(ir === 'b0000, "Assert 2688 : < ir !== 'b0000 >");	// Vector No: 672
verify(op === 'b00000000, "Assert 2689 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2690 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 2691 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 674
#2;

verify(ir === 'b1000, "Assert 2692 : < ir !== 'b1000 >");	// Vector No: 673
verify(op === 'b00000000, "Assert 2693 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2694 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2695 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 675
#2;

verify(ir === 'b0000, "Assert 2696 : < ir !== 'b0000 >");	// Vector No: 674
verify(op === 'b00000000, "Assert 2697 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2698 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 2699 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 676
#2;

verify(ir === 'b0000, "Assert 2700 : < ir !== 'b0000 >");	// Vector No: 675
verify(op === 'b00000000, "Assert 2701 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2702 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2703 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 677
#2;

verify(ir === 'b0000, "Assert 2704 : < ir !== 'b0000 >");	// Vector No: 676
verify(op === 'b00000000, "Assert 2705 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2706 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 2707 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 678
#2;

verify(ir === 'b1000, "Assert 2708 : < ir !== 'b1000 >");	// Vector No: 677
verify(op === 'b00000000, "Assert 2709 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2710 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2711 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 679
#2;

verify(ir === 'b0000, "Assert 2712 : < ir !== 'b0000 >");	// Vector No: 678
verify(op === 'b00000000, "Assert 2713 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2714 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 2715 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 680
#2;

verify(ir === 'b0000, "Assert 2716 : < ir !== 'b0000 >");	// Vector No: 679
verify(op === 'b00000000, "Assert 2717 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2718 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2719 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 681
#2;

verify(ir === 'b0000, "Assert 2720 : < ir !== 'b0000 >");	// Vector No: 680
verify(op === 'b00000000, "Assert 2721 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2722 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 2723 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 682
#2;

verify(ir === 'b1000, "Assert 2724 : < ir !== 'b1000 >");	// Vector No: 681
verify(op === 'b00000000, "Assert 2725 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2726 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2727 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 683
#2;

verify(ir === 'b0000, "Assert 2728 : < ir !== 'b0000 >");	// Vector No: 682
verify(op === 'b00000000, "Assert 2729 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2730 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 2731 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 684
#2;

verify(ir === 'b0000, "Assert 2732 : < ir !== 'b0000 >");	// Vector No: 683
verify(op === 'b00000000, "Assert 2733 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2734 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2735 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 685
#2;

verify(ir === 'b0000, "Assert 2736 : < ir !== 'b0000 >");	// Vector No: 684
verify(op === 'b00000000, "Assert 2737 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2738 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 2739 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 686
#2;

verify(ir === 'b1000, "Assert 2740 : < ir !== 'b1000 >");	// Vector No: 685
verify(op === 'b00000000, "Assert 2741 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2742 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2743 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 687
#2;

verify(ir === 'b0000, "Assert 2744 : < ir !== 'b0000 >");	// Vector No: 686
verify(op === 'b00000000, "Assert 2745 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2746 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 2747 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 688
#2;

verify(ir === 'b0000, "Assert 2748 : < ir !== 'b0000 >");	// Vector No: 687
verify(op === 'b00000000, "Assert 2749 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2750 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2751 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 689
#2;

verify(ir === 'b0000, "Assert 2752 : < ir !== 'b0000 >");	// Vector No: 688
verify(op === 'b00000000, "Assert 2753 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2754 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 2755 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 690
#2;

verify(ir === 'b1000, "Assert 2756 : < ir !== 'b1000 >");	// Vector No: 689
verify(op === 'b00000000, "Assert 2757 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2758 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2759 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 691
#2;

verify(ir === 'b0000, "Assert 2760 : < ir !== 'b0000 >");	// Vector No: 690
verify(op === 'b00000000, "Assert 2761 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2762 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 2763 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 692
#2;

verify(ir === 'b0000, "Assert 2764 : < ir !== 'b0000 >");	// Vector No: 691
verify(op === 'b00000000, "Assert 2765 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2766 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2767 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 693
#2;

verify(ir === 'b0000, "Assert 2768 : < ir !== 'b0000 >");	// Vector No: 692
verify(op === 'b00000000, "Assert 2769 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2770 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 2771 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 694
#2;

verify(ir === 'b1000, "Assert 2772 : < ir !== 'b1000 >");	// Vector No: 693
verify(op === 'b00000000, "Assert 2773 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2774 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2775 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 695
#2;

verify(ir === 'b0000, "Assert 2776 : < ir !== 'b0000 >");	// Vector No: 694
verify(op === 'b00000000, "Assert 2777 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2778 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 2779 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 696
#2;

verify(ir === 'b0000, "Assert 2780 : < ir !== 'b0000 >");	// Vector No: 695
verify(op === 'b00000000, "Assert 2781 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2782 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2783 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 697
#2;

verify(ir === 'b0000, "Assert 2784 : < ir !== 'b0000 >");	// Vector No: 696
verify(op === 'b00000000, "Assert 2785 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2786 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 2787 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 698
#2;

verify(ir === 'b1000, "Assert 2788 : < ir !== 'b1000 >");	// Vector No: 697
verify(op === 'b00000000, "Assert 2789 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2790 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2791 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 699
#2;

verify(ir === 'b0000, "Assert 2792 : < ir !== 'b0000 >");	// Vector No: 698
verify(op === 'b00000000, "Assert 2793 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2794 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 2795 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 700
#2;

verify(ir === 'b0000, "Assert 2796 : < ir !== 'b0000 >");	// Vector No: 699
verify(op === 'b00000000, "Assert 2797 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2798 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2799 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 701
#2;

verify(ir === 'b0000, "Assert 2800 : < ir !== 'b0000 >");	// Vector No: 700
verify(op === 'b00000000, "Assert 2801 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2802 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 2803 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 702
#2;

verify(ir === 'b1000, "Assert 2804 : < ir !== 'b1000 >");	// Vector No: 701
verify(op === 'b00000000, "Assert 2805 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2806 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2807 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000010000000000000000000000000000000:1:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 703
#2;

verify(ir === 'b0000, "Assert 2808 : < ir !== 'b0000 >");	// Vector No: 702
verify(op === 'b00000001, "Assert 2809 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 2810 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2811 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 704
#2;

verify(ir === 'b0000, "Assert 2812 : < ir !== 'b0000 >");	// Vector No: 703
verify(op === 'b00000000, "Assert 2813 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2814 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2815 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000010000000000000000000000000000000:0:0:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 705
#2;

verify(ir === 'b0000, "Assert 2816 : < ir !== 'b0000 >");	// Vector No: 704
verify(op === 'b00000000, "Assert 2817 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2818 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 2819 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 706
#2;

verify(ir === 'b1000, "Assert 2820 : < ir !== 'b1000 >");	// Vector No: 705
verify(op === 'b00000000, "Assert 2821 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2822 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2823 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000010000000000000000000000000000000:1:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 707
#2;

verify(ir === 'b0000, "Assert 2824 : < ir !== 'b0000 >");	// Vector No: 706
verify(op === 'b00000010, "Assert 2825 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 2826 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2827 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 708
#2;

verify(ir === 'b0000, "Assert 2828 : < ir !== 'b0000 >");	// Vector No: 707
verify(op === 'b00000000, "Assert 2829 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2830 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2831 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000010000000000000000000000000000000:0:0:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 709
#2;

verify(ir === 'b0000, "Assert 2832 : < ir !== 'b0000 >");	// Vector No: 708
verify(op === 'b00000000, "Assert 2833 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2834 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 2835 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 710
#2;

verify(ir === 'b1000, "Assert 2836 : < ir !== 'b1000 >");	// Vector No: 709
verify(op === 'b00000000, "Assert 2837 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2838 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2839 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000010000000000000000000000000000000:1:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 711
#2;

verify(ir === 'b0000, "Assert 2840 : < ir !== 'b0000 >");	// Vector No: 710
verify(op === 'b00000100, "Assert 2841 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 2842 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2843 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 712
#2;

verify(ir === 'b0000, "Assert 2844 : < ir !== 'b0000 >");	// Vector No: 711
verify(op === 'b00000000, "Assert 2845 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2846 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2847 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000010000000000000000000000000000000:0:0:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 713
#2;

verify(ir === 'b0000, "Assert 2848 : < ir !== 'b0000 >");	// Vector No: 712
verify(op === 'b00000000, "Assert 2849 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2850 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 2851 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 714
#2;

verify(ir === 'b1000, "Assert 2852 : < ir !== 'b1000 >");	// Vector No: 713
verify(op === 'b00000000, "Assert 2853 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2854 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2855 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000010000000000000000000000000000000:1:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 715
#2;

verify(ir === 'b0000, "Assert 2856 : < ir !== 'b0000 >");	// Vector No: 714
verify(op === 'b00001000, "Assert 2857 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 2858 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2859 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 716
#2;

verify(ir === 'b0000, "Assert 2860 : < ir !== 'b0000 >");	// Vector No: 715
verify(op === 'b00000000, "Assert 2861 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2862 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2863 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000010000000000000000000000000000000:0:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 717
#2;

verify(ir === 'b0000, "Assert 2864 : < ir !== 'b0000 >");	// Vector No: 716
verify(op === 'b00000001, "Assert 2865 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 2866 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2867 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 718
#2;

verify(ir === 'b1000, "Assert 2868 : < ir !== 'b1000 >");	// Vector No: 717
verify(op === 'b00000000, "Assert 2869 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2870 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2871 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000010000000000000000000000000000000:1:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 719
#2;

verify(ir === 'b0000, "Assert 2872 : < ir !== 'b0000 >");	// Vector No: 718
verify(op === 'b00010000, "Assert 2873 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 2874 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2875 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 720
#2;

verify(ir === 'b0000, "Assert 2876 : < ir !== 'b0000 >");	// Vector No: 719
verify(op === 'b00000000, "Assert 2877 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2878 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2879 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000010000000000000000000000000000000:0:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 721
#2;

verify(ir === 'b0000, "Assert 2880 : < ir !== 'b0000 >");	// Vector No: 720
verify(op === 'b00000010, "Assert 2881 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 2882 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2883 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 722
#2;

verify(ir === 'b1000, "Assert 2884 : < ir !== 'b1000 >");	// Vector No: 721
verify(op === 'b00000000, "Assert 2885 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2886 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2887 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000010000000000000000000000000000000:1:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 723
#2;

verify(ir === 'b0000, "Assert 2888 : < ir !== 'b0000 >");	// Vector No: 722
verify(op === 'b00100000, "Assert 2889 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 2890 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2891 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 724
#2;

verify(ir === 'b0000, "Assert 2892 : < ir !== 'b0000 >");	// Vector No: 723
verify(op === 'b00000000, "Assert 2893 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2894 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2895 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000010000000000000000000000000000000:0:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 725
#2;

verify(ir === 'b0000, "Assert 2896 : < ir !== 'b0000 >");	// Vector No: 724
verify(op === 'b00000100, "Assert 2897 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 2898 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2899 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 726
#2;

verify(ir === 'b1000, "Assert 2900 : < ir !== 'b1000 >");	// Vector No: 725
verify(op === 'b00000000, "Assert 2901 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2902 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2903 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000010000000000000000000000000000000:1:0:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 727
#2;

verify(ir === 'b0000, "Assert 2904 : < ir !== 'b0000 >");	// Vector No: 726
verify(op === 'b01000000, "Assert 2905 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 2906 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 2907 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 728
#2;

verify(ir === 'b0000, "Assert 2908 : < ir !== 'b0000 >");	// Vector No: 727
verify(op === 'b00000000, "Assert 2909 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2910 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2911 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000010000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 729
#2;

verify(ir === 'b0000, "Assert 2912 : < ir !== 'b0000 >");	// Vector No: 728
verify(op === 'b00001000, "Assert 2913 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 2914 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2915 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 730
#2;

verify(ir === 'b1000, "Assert 2916 : < ir !== 'b1000 >");	// Vector No: 729
verify(op === 'b00000000, "Assert 2917 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2918 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2919 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000010000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 731
#2;

verify(ir === 'b0000, "Assert 2920 : < ir !== 'b0000 >");	// Vector No: 730
verify(op === 'b10000000, "Assert 2921 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 2922 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2923 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 732
#2;

verify(ir === 'b0000, "Assert 2924 : < ir !== 'b0000 >");	// Vector No: 731
verify(op === 'b00000000, "Assert 2925 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2926 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2927 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000010000000000000000000000000000000:0:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 733
#2;

verify(ir === 'b0000, "Assert 2928 : < ir !== 'b0000 >");	// Vector No: 732
verify(op === 'b00010000, "Assert 2929 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 2930 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2931 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 734
#2;

verify(ir === 'b1000, "Assert 2932 : < ir !== 'b1000 >");	// Vector No: 733
verify(op === 'b00000000, "Assert 2933 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2934 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2935 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000010000000000000000000000000000000:1:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 735
#2;

verify(ir === 'b0001, "Assert 2936 : < ir !== 'b0001 >");	// Vector No: 734
verify(op === 'b00000000, "Assert 2937 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2938 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2939 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 736
#2;

verify(ir === 'b0000, "Assert 2940 : < ir !== 'b0000 >");	// Vector No: 735
verify(op === 'b00000000, "Assert 2941 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2942 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2943 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000010000000000000000000000000000000:0:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 737
#2;

verify(ir === 'b0000, "Assert 2944 : < ir !== 'b0000 >");	// Vector No: 736
verify(op === 'b00100000, "Assert 2945 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 2946 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2947 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 738
#2;

verify(ir === 'b1000, "Assert 2948 : < ir !== 'b1000 >");	// Vector No: 737
verify(op === 'b00000000, "Assert 2949 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2950 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2951 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000010000000000000000000000000000000:1:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 739
#2;

verify(ir === 'b0010, "Assert 2952 : < ir !== 'b0010 >");	// Vector No: 738
verify(op === 'b00000000, "Assert 2953 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2954 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2955 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 740
#2;

verify(ir === 'b0000, "Assert 2956 : < ir !== 'b0000 >");	// Vector No: 739
verify(op === 'b00000000, "Assert 2957 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2958 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2959 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000010000000000000000000000000000000:0:0:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 741
#2;

verify(ir === 'b0000, "Assert 2960 : < ir !== 'b0000 >");	// Vector No: 740
verify(op === 'b01000000, "Assert 2961 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 2962 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2963 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 742
#2;

verify(ir === 'b1000, "Assert 2964 : < ir !== 'b1000 >");	// Vector No: 741
verify(op === 'b00000000, "Assert 2965 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2966 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2967 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000010000000000000000000000000000000:1:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 743
#2;

verify(ir === 'b0100, "Assert 2968 : < ir !== 'b0100 >");	// Vector No: 742
verify(op === 'b00000000, "Assert 2969 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2970 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2971 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 744
#2;

verify(ir === 'b0000, "Assert 2972 : < ir !== 'b0000 >");	// Vector No: 743
verify(op === 'b00000000, "Assert 2973 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2974 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2975 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000010000000000000000000000000000000:0:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 745
#2;

verify(ir === 'b0000, "Assert 2976 : < ir !== 'b0000 >");	// Vector No: 744
verify(op === 'b10000000, "Assert 2977 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 2978 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2979 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 746
#2;

verify(ir === 'b1000, "Assert 2980 : < ir !== 'b1000 >");	// Vector No: 745
verify(op === 'b00000000, "Assert 2981 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2982 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2983 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 747
#2;

verify(ir === 'b0000, "Assert 2984 : < ir !== 'b0000 >");	// Vector No: 746
verify(op === 'b00000000, "Assert 2985 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2986 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2987 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 748
#2;

verify(ir === 'b0000, "Assert 2988 : < ir !== 'b0000 >");	// Vector No: 747
verify(op === 'b00000000, "Assert 2989 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2990 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2991 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000010000000000000000000000000000000:0:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 749
#2;

verify(ir === 'b0001, "Assert 2992 : < ir !== 'b0001 >");	// Vector No: 748
verify(op === 'b00000000, "Assert 2993 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2994 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2995 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 750
#2;

verify(ir === 'b1000, "Assert 2996 : < ir !== 'b1000 >");	// Vector No: 749
verify(op === 'b00000000, "Assert 2997 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 2998 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 2999 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 751
#2;

verify(ir === 'b0000, "Assert 3000 : < ir !== 'b0000 >");	// Vector No: 750
verify(op === 'b00000000, "Assert 3001 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3002 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3003 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 752
#2;

verify(ir === 'b0000, "Assert 3004 : < ir !== 'b0000 >");	// Vector No: 751
verify(op === 'b00000000, "Assert 3005 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3006 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3007 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000010000000000000000000000000000000:0:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 753
#2;

verify(ir === 'b0010, "Assert 3008 : < ir !== 'b0010 >");	// Vector No: 752
verify(op === 'b00000000, "Assert 3009 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3010 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3011 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 754
#2;

verify(ir === 'b1000, "Assert 3012 : < ir !== 'b1000 >");	// Vector No: 753
verify(op === 'b00000000, "Assert 3013 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3014 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3015 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 755
#2;

verify(ir === 'b0000, "Assert 3016 : < ir !== 'b0000 >");	// Vector No: 754
verify(op === 'b00000000, "Assert 3017 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3018 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3019 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 756
#2;

verify(ir === 'b0000, "Assert 3020 : < ir !== 'b0000 >");	// Vector No: 755
verify(op === 'b00000000, "Assert 3021 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3022 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3023 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000010000000000000000000000000000000:0:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 757
#2;

verify(ir === 'b0100, "Assert 3024 : < ir !== 'b0100 >");	// Vector No: 756
verify(op === 'b00000000, "Assert 3025 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3026 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3027 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 758
#2;

verify(ir === 'b1000, "Assert 3028 : < ir !== 'b1000 >");	// Vector No: 757
verify(op === 'b00000000, "Assert 3029 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3030 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3031 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000010000000000000000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 759
#2;

verify(ir === 'b0000, "Assert 3032 : < ir !== 'b0000 >");	// Vector No: 758
verify(op === 'b00000000, "Assert 3033 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3034 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3035 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 760
#2;

verify(ir === 'b0000, "Assert 3036 : < ir !== 'b0000 >");	// Vector No: 759
verify(op === 'b00000000, "Assert 3037 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3038 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3039 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000010000000000000000000000000000000:0:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 761
#2;

verify(ir === 'b1000, "Assert 3040 : < ir !== 'b1000 >");	// Vector No: 760
verify(op === 'b00000000, "Assert 3041 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3042 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3043 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 762
#2;

verify(ir === 'b1000, "Assert 3044 : < ir !== 'b1000 >");	// Vector No: 761
verify(op === 'b00000000, "Assert 3045 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3046 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3047 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000010000000000000000000000000000000:1:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 763
#2;

verify(ir === 'b1000, "Assert 3048 : < ir !== 'b1000 >");	// Vector No: 762
verify(op === 'b00000000, "Assert 3049 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3050 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3051 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 764
#2;

verify(ir === 'b0000, "Assert 3052 : < ir !== 'b0000 >");	// Vector No: 763
verify(op === 'b00000000, "Assert 3053 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3054 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3055 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000001:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 765
#2;

verify(ir === 'b0000, "Assert 3056 : < ir !== 'b0000 >");	// Vector No: 764
verify(op === 'b00001000, "Assert 3057 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3058 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3059 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000001:0:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 766
#2;

verify(ir === 'b0000, "Assert 3060 : < ir !== 'b0000 >");	// Vector No: 765
verify(op === 'b00000000, "Assert 3061 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3062 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 3063 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000001:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 767
#2;

verify(ir === 'b0000, "Assert 3064 : < ir !== 'b0000 >");	// Vector No: 766
verify(op === 'b10000000, "Assert 3065 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3066 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3067 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000001:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 768
#2;

verify(ir === 'b0000, "Assert 3068 : < ir !== 'b0000 >");	// Vector No: 767
verify(op === 'b00000000, "Assert 3069 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3070 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3071 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000010:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 769
#2;

verify(ir === 'b0000, "Assert 3072 : < ir !== 'b0000 >");	// Vector No: 768
verify(op === 'b00001000, "Assert 3073 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3074 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3075 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000010:0:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 770
#2;

verify(ir === 'b0000, "Assert 3076 : < ir !== 'b0000 >");	// Vector No: 769
verify(op === 'b00000000, "Assert 3077 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3078 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 3079 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000010:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 771
#2;

verify(ir === 'b0000, "Assert 3080 : < ir !== 'b0000 >");	// Vector No: 770
verify(op === 'b10000000, "Assert 3081 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3082 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3083 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000010:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 772
#2;

verify(ir === 'b0000, "Assert 3084 : < ir !== 'b0000 >");	// Vector No: 771
verify(op === 'b00000000, "Assert 3085 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3086 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3087 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000100:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 773
#2;

verify(ir === 'b0000, "Assert 3088 : < ir !== 'b0000 >");	// Vector No: 772
verify(op === 'b00001000, "Assert 3089 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3090 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3091 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000100:0:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 774
#2;

verify(ir === 'b0000, "Assert 3092 : < ir !== 'b0000 >");	// Vector No: 773
verify(op === 'b00000000, "Assert 3093 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3094 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 3095 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000100:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 775
#2;

verify(ir === 'b0000, "Assert 3096 : < ir !== 'b0000 >");	// Vector No: 774
verify(op === 'b10000000, "Assert 3097 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3098 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3099 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000000100:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 776
#2;

verify(ir === 'b0000, "Assert 3100 : < ir !== 'b0000 >");	// Vector No: 775
verify(op === 'b00000000, "Assert 3101 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3102 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3103 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000001000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 777
#2;

verify(ir === 'b0000, "Assert 3104 : < ir !== 'b0000 >");	// Vector No: 776
verify(op === 'b00001000, "Assert 3105 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3106 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3107 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000001000:0:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 778
#2;

verify(ir === 'b0000, "Assert 3108 : < ir !== 'b0000 >");	// Vector No: 777
verify(op === 'b00000000, "Assert 3109 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3110 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 3111 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000001000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 779
#2;

verify(ir === 'b0000, "Assert 3112 : < ir !== 'b0000 >");	// Vector No: 778
verify(op === 'b10000000, "Assert 3113 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3114 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3115 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000001000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 780
#2;

verify(ir === 'b0000, "Assert 3116 : < ir !== 'b0000 >");	// Vector No: 779
verify(op === 'b00000000, "Assert 3117 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3118 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3119 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000010000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 781
#2;

verify(ir === 'b0000, "Assert 3120 : < ir !== 'b0000 >");	// Vector No: 780
verify(op === 'b00001000, "Assert 3121 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3122 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3123 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000010000:0:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 782
#2;

verify(ir === 'b0000, "Assert 3124 : < ir !== 'b0000 >");	// Vector No: 781
verify(op === 'b00000000, "Assert 3125 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3126 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 3127 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000010000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 783
#2;

verify(ir === 'b0000, "Assert 3128 : < ir !== 'b0000 >");	// Vector No: 782
verify(op === 'b10000000, "Assert 3129 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3130 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3131 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000010000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 784
#2;

verify(ir === 'b0000, "Assert 3132 : < ir !== 'b0000 >");	// Vector No: 783
verify(op === 'b00000000, "Assert 3133 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3134 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3135 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000100000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 785
#2;

verify(ir === 'b0000, "Assert 3136 : < ir !== 'b0000 >");	// Vector No: 784
verify(op === 'b00001000, "Assert 3137 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3138 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3139 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000100000:0:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 786
#2;

verify(ir === 'b0000, "Assert 3140 : < ir !== 'b0000 >");	// Vector No: 785
verify(op === 'b00000000, "Assert 3141 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3142 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 3143 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000100000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 787
#2;

verify(ir === 'b0000, "Assert 3144 : < ir !== 'b0000 >");	// Vector No: 786
verify(op === 'b10000000, "Assert 3145 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3146 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3147 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000000100000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 788
#2;

verify(ir === 'b0000, "Assert 3148 : < ir !== 'b0000 >");	// Vector No: 787
verify(op === 'b00000000, "Assert 3149 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3150 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3151 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000001000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 789
#2;

verify(ir === 'b0000, "Assert 3152 : < ir !== 'b0000 >");	// Vector No: 788
verify(op === 'b00001000, "Assert 3153 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3154 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3155 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000001000000:0:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 790
#2;

verify(ir === 'b0000, "Assert 3156 : < ir !== 'b0000 >");	// Vector No: 789
verify(op === 'b00000000, "Assert 3157 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3158 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 3159 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000001000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 791
#2;

verify(ir === 'b0000, "Assert 3160 : < ir !== 'b0000 >");	// Vector No: 790
verify(op === 'b10000000, "Assert 3161 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3162 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3163 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000001000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 792
#2;

verify(ir === 'b0000, "Assert 3164 : < ir !== 'b0000 >");	// Vector No: 791
verify(op === 'b00000000, "Assert 3165 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3166 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3167 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000010000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 793
#2;

verify(ir === 'b0000, "Assert 3168 : < ir !== 'b0000 >");	// Vector No: 792
verify(op === 'b00001000, "Assert 3169 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3170 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3171 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000010000000:0:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 794
#2;

verify(ir === 'b0000, "Assert 3172 : < ir !== 'b0000 >");	// Vector No: 793
verify(op === 'b00000000, "Assert 3173 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3174 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 3175 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000010000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 795
#2;

verify(ir === 'b0000, "Assert 3176 : < ir !== 'b0000 >");	// Vector No: 794
verify(op === 'b10000000, "Assert 3177 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3178 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3179 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000010000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 796
#2;

verify(ir === 'b0000, "Assert 3180 : < ir !== 'b0000 >");	// Vector No: 795
verify(op === 'b00000000, "Assert 3181 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3182 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3183 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000100000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 797
#2;

verify(ir === 'b0000, "Assert 3184 : < ir !== 'b0000 >");	// Vector No: 796
verify(op === 'b00001000, "Assert 3185 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3186 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3187 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000100000000:0:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 798
#2;

verify(ir === 'b0000, "Assert 3188 : < ir !== 'b0000 >");	// Vector No: 797
verify(op === 'b00000000, "Assert 3189 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3190 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 3191 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000100000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 799
#2;

verify(ir === 'b0000, "Assert 3192 : < ir !== 'b0000 >");	// Vector No: 798
verify(op === 'b10000000, "Assert 3193 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3194 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3195 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000000100000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 800
#2;

verify(ir === 'b0000, "Assert 3196 : < ir !== 'b0000 >");	// Vector No: 799
verify(op === 'b00000000, "Assert 3197 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3198 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3199 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000001000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 801
#2;

verify(ir === 'b0000, "Assert 3200 : < ir !== 'b0000 >");	// Vector No: 800
verify(op === 'b00001000, "Assert 3201 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3202 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3203 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000001000000000:0:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 802
#2;

verify(ir === 'b0000, "Assert 3204 : < ir !== 'b0000 >");	// Vector No: 801
verify(op === 'b00000000, "Assert 3205 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3206 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 3207 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000001000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 803
#2;

verify(ir === 'b0000, "Assert 3208 : < ir !== 'b0000 >");	// Vector No: 802
verify(op === 'b10000000, "Assert 3209 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3210 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3211 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000001000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 804
#2;

verify(ir === 'b0000, "Assert 3212 : < ir !== 'b0000 >");	// Vector No: 803
verify(op === 'b00000000, "Assert 3213 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3214 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3215 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000010000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 805
#2;

verify(ir === 'b0000, "Assert 3216 : < ir !== 'b0000 >");	// Vector No: 804
verify(op === 'b00001000, "Assert 3217 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3218 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3219 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000010000000000:0:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 806
#2;

verify(ir === 'b0000, "Assert 3220 : < ir !== 'b0000 >");	// Vector No: 805
verify(op === 'b00000000, "Assert 3221 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3222 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 3223 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000010000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 807
#2;

verify(ir === 'b0000, "Assert 3224 : < ir !== 'b0000 >");	// Vector No: 806
verify(op === 'b10000000, "Assert 3225 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3226 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3227 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000010000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 808
#2;

verify(ir === 'b0000, "Assert 3228 : < ir !== 'b0000 >");	// Vector No: 807
verify(op === 'b00000000, "Assert 3229 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3230 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3231 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000100000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 809
#2;

verify(ir === 'b0000, "Assert 3232 : < ir !== 'b0000 >");	// Vector No: 808
verify(op === 'b00001000, "Assert 3233 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3234 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3235 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000100000000000:0:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 810
#2;

verify(ir === 'b0000, "Assert 3236 : < ir !== 'b0000 >");	// Vector No: 809
verify(op === 'b00000000, "Assert 3237 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3238 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 3239 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000100000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 811
#2;

verify(ir === 'b0000, "Assert 3240 : < ir !== 'b0000 >");	// Vector No: 810
verify(op === 'b10000000, "Assert 3241 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3242 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3243 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000000100000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 812
#2;

verify(ir === 'b0000, "Assert 3244 : < ir !== 'b0000 >");	// Vector No: 811
verify(op === 'b00000000, "Assert 3245 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3246 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3247 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000001000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 813
#2;

verify(ir === 'b0000, "Assert 3248 : < ir !== 'b0000 >");	// Vector No: 812
verify(op === 'b00001000, "Assert 3249 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3250 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3251 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000001000000000000:0:1:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 814
#2;

verify(ir === 'b0000, "Assert 3252 : < ir !== 'b0000 >");	// Vector No: 813
verify(op === 'b00000000, "Assert 3253 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3254 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 3255 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000001000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 815
#2;

verify(ir === 'b0000, "Assert 3256 : < ir !== 'b0000 >");	// Vector No: 814
verify(op === 'b10000000, "Assert 3257 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3258 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3259 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000001000000000000:1:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 816
#2;

verify(ir === 'b0000, "Assert 3260 : < ir !== 'b0000 >");	// Vector No: 815
verify(op === 'b00000000, "Assert 3261 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3262 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 3263 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000010000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 817
#2;

verify(ir === 'b0000, "Assert 3264 : < ir !== 'b0000 >");	// Vector No: 816
verify(op === 'b00001000, "Assert 3265 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3266 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3267 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000010000000000000:0:1:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 818
#2;

verify(ir === 'b0000, "Assert 3268 : < ir !== 'b0000 >");	// Vector No: 817
verify(op === 'b00000000, "Assert 3269 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3270 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 3271 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000010000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 819
#2;

verify(ir === 'b0000, "Assert 3272 : < ir !== 'b0000 >");	// Vector No: 818
verify(op === 'b10000000, "Assert 3273 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3274 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3275 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000010000000000000:1:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 820
#2;

verify(ir === 'b0000, "Assert 3276 : < ir !== 'b0000 >");	// Vector No: 819
verify(op === 'b00000000, "Assert 3277 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3278 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 3279 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000100000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 821
#2;

verify(ir === 'b0000, "Assert 3280 : < ir !== 'b0000 >");	// Vector No: 820
verify(op === 'b00001000, "Assert 3281 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3282 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3283 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000100000000000000:0:1:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 822
#2;

verify(ir === 'b0000, "Assert 3284 : < ir !== 'b0000 >");	// Vector No: 821
verify(op === 'b00000000, "Assert 3285 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3286 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 3287 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000100000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 823
#2;

verify(ir === 'b0000, "Assert 3288 : < ir !== 'b0000 >");	// Vector No: 822
verify(op === 'b10000000, "Assert 3289 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3290 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3291 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000000100000000000000:1:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 824
#2;

verify(ir === 'b0000, "Assert 3292 : < ir !== 'b0000 >");	// Vector No: 823
verify(op === 'b00000000, "Assert 3293 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3294 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 3295 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000001000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 825
#2;

verify(ir === 'b0000, "Assert 3296 : < ir !== 'b0000 >");	// Vector No: 824
verify(op === 'b00001000, "Assert 3297 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3298 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3299 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000001000000000000000:0:1:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 826
#2;

verify(ir === 'b0000, "Assert 3300 : < ir !== 'b0000 >");	// Vector No: 825
verify(op === 'b00000000, "Assert 3301 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3302 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 3303 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000001000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 827
#2;

verify(ir === 'b0000, "Assert 3304 : < ir !== 'b0000 >");	// Vector No: 826
verify(op === 'b10000000, "Assert 3305 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3306 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3307 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000001000000000000000:1:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 828
#2;

verify(ir === 'b0000, "Assert 3308 : < ir !== 'b0000 >");	// Vector No: 827
verify(op === 'b00000000, "Assert 3309 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3310 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 3311 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000010000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 829
#2;

verify(ir === 'b0000, "Assert 3312 : < ir !== 'b0000 >");	// Vector No: 828
verify(op === 'b00001000, "Assert 3313 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3314 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3315 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000010000000000000000:0:1:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 830
#2;

verify(ir === 'b0000, "Assert 3316 : < ir !== 'b0000 >");	// Vector No: 829
verify(op === 'b00000000, "Assert 3317 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3318 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 3319 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000010000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 831
#2;

verify(ir === 'b0000, "Assert 3320 : < ir !== 'b0000 >");	// Vector No: 830
verify(op === 'b10000000, "Assert 3321 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3322 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3323 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000010000000000000000:1:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 832
#2;

verify(ir === 'b0000, "Assert 3324 : < ir !== 'b0000 >");	// Vector No: 831
verify(op === 'b00000000, "Assert 3325 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3326 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 3327 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000100000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 833
#2;

verify(ir === 'b0000, "Assert 3328 : < ir !== 'b0000 >");	// Vector No: 832
verify(op === 'b00001000, "Assert 3329 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3330 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3331 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000100000000000000000:0:1:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 834
#2;

verify(ir === 'b0000, "Assert 3332 : < ir !== 'b0000 >");	// Vector No: 833
verify(op === 'b00000000, "Assert 3333 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3334 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 3335 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000100000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 835
#2;

verify(ir === 'b0000, "Assert 3336 : < ir !== 'b0000 >");	// Vector No: 834
verify(op === 'b10000000, "Assert 3337 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3338 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3339 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000000100000000000000000:1:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 836
#2;

verify(ir === 'b0000, "Assert 3340 : < ir !== 'b0000 >");	// Vector No: 835
verify(op === 'b00000000, "Assert 3341 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3342 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 3343 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000001000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 837
#2;

verify(ir === 'b0000, "Assert 3344 : < ir !== 'b0000 >");	// Vector No: 836
verify(op === 'b00001000, "Assert 3345 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3346 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3347 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000001000000000000000000:0:1:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 838
#2;

verify(ir === 'b0000, "Assert 3348 : < ir !== 'b0000 >");	// Vector No: 837
verify(op === 'b00000000, "Assert 3349 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3350 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 3351 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000001000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 839
#2;

verify(ir === 'b0000, "Assert 3352 : < ir !== 'b0000 >");	// Vector No: 838
verify(op === 'b10000000, "Assert 3353 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3354 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3355 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000001000000000000000000:1:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 840
#2;

verify(ir === 'b0000, "Assert 3356 : < ir !== 'b0000 >");	// Vector No: 839
verify(op === 'b00000000, "Assert 3357 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3358 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 3359 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000010000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 841
#2;

verify(ir === 'b0000, "Assert 3360 : < ir !== 'b0000 >");	// Vector No: 840
verify(op === 'b00001000, "Assert 3361 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3362 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3363 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000010000000000000000000:0:1:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 842
#2;

verify(ir === 'b0000, "Assert 3364 : < ir !== 'b0000 >");	// Vector No: 841
verify(op === 'b00000000, "Assert 3365 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3366 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 3367 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000010000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 843
#2;

verify(ir === 'b0000, "Assert 3368 : < ir !== 'b0000 >");	// Vector No: 842
verify(op === 'b10000000, "Assert 3369 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3370 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3371 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000010000000000000000000:1:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 844
#2;

verify(ir === 'b0000, "Assert 3372 : < ir !== 'b0000 >");	// Vector No: 843
verify(op === 'b00000000, "Assert 3373 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3374 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 3375 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000100000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 845
#2;

verify(ir === 'b0000, "Assert 3376 : < ir !== 'b0000 >");	// Vector No: 844
verify(op === 'b00001000, "Assert 3377 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3378 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3379 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000100000000000000000000:0:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 846
#2;

verify(ir === 'b0000, "Assert 3380 : < ir !== 'b0000 >");	// Vector No: 845
verify(op === 'b00000001, "Assert 3381 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 3382 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3383 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000100000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 847
#2;

verify(ir === 'b0000, "Assert 3384 : < ir !== 'b0000 >");	// Vector No: 846
verify(op === 'b10000000, "Assert 3385 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3386 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3387 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000000100000000000000000000:1:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 848
#2;

verify(ir === 'b0000, "Assert 3388 : < ir !== 'b0000 >");	// Vector No: 847
verify(op === 'b00000000, "Assert 3389 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3390 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 3391 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000001000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 849
#2;

verify(ir === 'b0000, "Assert 3392 : < ir !== 'b0000 >");	// Vector No: 848
verify(op === 'b00001000, "Assert 3393 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3394 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3395 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000001000000000000000000000:0:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 850
#2;

verify(ir === 'b0000, "Assert 3396 : < ir !== 'b0000 >");	// Vector No: 849
verify(op === 'b00000010, "Assert 3397 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 3398 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3399 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000001000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 851
#2;

verify(ir === 'b0000, "Assert 3400 : < ir !== 'b0000 >");	// Vector No: 850
verify(op === 'b10000000, "Assert 3401 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3402 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3403 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000001000000000000000000000:1:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 852
#2;

verify(ir === 'b0000, "Assert 3404 : < ir !== 'b0000 >");	// Vector No: 851
verify(op === 'b00000000, "Assert 3405 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3406 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 3407 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000010000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 853
#2;

verify(ir === 'b0000, "Assert 3408 : < ir !== 'b0000 >");	// Vector No: 852
verify(op === 'b00001000, "Assert 3409 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3410 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3411 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000010000000000000000000000:0:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 854
#2;

verify(ir === 'b0000, "Assert 3412 : < ir !== 'b0000 >");	// Vector No: 853
verify(op === 'b00000100, "Assert 3413 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 3414 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3415 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000010000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 855
#2;

verify(ir === 'b0000, "Assert 3416 : < ir !== 'b0000 >");	// Vector No: 854
verify(op === 'b10000000, "Assert 3417 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3418 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3419 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000010000000000000000000000:1:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 856
#2;

verify(ir === 'b0000, "Assert 3420 : < ir !== 'b0000 >");	// Vector No: 855
verify(op === 'b00000000, "Assert 3421 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3422 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 3423 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000100000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 857
#2;

verify(ir === 'b0000, "Assert 3424 : < ir !== 'b0000 >");	// Vector No: 856
verify(op === 'b00001000, "Assert 3425 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3426 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3427 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000100000000000000000000000:0:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 858
#2;

verify(ir === 'b0000, "Assert 3428 : < ir !== 'b0000 >");	// Vector No: 857
verify(op === 'b00001000, "Assert 3429 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3430 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3431 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000100000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 859
#2;

verify(ir === 'b0000, "Assert 3432 : < ir !== 'b0000 >");	// Vector No: 858
verify(op === 'b10000000, "Assert 3433 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3434 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3435 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000000100000000000000000000000:1:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 860
#2;

verify(ir === 'b0000, "Assert 3436 : < ir !== 'b0000 >");	// Vector No: 859
verify(op === 'b00000000, "Assert 3437 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3438 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 3439 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000001000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 861
#2;

verify(ir === 'b0000, "Assert 3440 : < ir !== 'b0000 >");	// Vector No: 860
verify(op === 'b00001000, "Assert 3441 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3442 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3443 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000001000000000000000000000000:0:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 862
#2;

verify(ir === 'b0000, "Assert 3444 : < ir !== 'b0000 >");	// Vector No: 861
verify(op === 'b00010000, "Assert 3445 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 3446 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3447 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000001000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 863
#2;

verify(ir === 'b0000, "Assert 3448 : < ir !== 'b0000 >");	// Vector No: 862
verify(op === 'b10000000, "Assert 3449 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3450 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3451 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000001000000000000000000000000:1:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 864
#2;

verify(ir === 'b0000, "Assert 3452 : < ir !== 'b0000 >");	// Vector No: 863
verify(op === 'b00000001, "Assert 3453 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 3454 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3455 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000010000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 865
#2;

verify(ir === 'b0000, "Assert 3456 : < ir !== 'b0000 >");	// Vector No: 864
verify(op === 'b00001000, "Assert 3457 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3458 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3459 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000010000000000000000000000000:0:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 866
#2;

verify(ir === 'b0000, "Assert 3460 : < ir !== 'b0000 >");	// Vector No: 865
verify(op === 'b00100000, "Assert 3461 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 3462 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3463 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000010000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 867
#2;

verify(ir === 'b0000, "Assert 3464 : < ir !== 'b0000 >");	// Vector No: 866
verify(op === 'b10000000, "Assert 3465 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3466 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3467 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000010000000000000000000000000:1:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 868
#2;

verify(ir === 'b0000, "Assert 3468 : < ir !== 'b0000 >");	// Vector No: 867
verify(op === 'b00000010, "Assert 3469 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 3470 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3471 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000100000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 869
#2;

verify(ir === 'b0000, "Assert 3472 : < ir !== 'b0000 >");	// Vector No: 868
verify(op === 'b00001000, "Assert 3473 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3474 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3475 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000100000000000000000000000000:0:1:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 870
#2;

verify(ir === 'b0000, "Assert 3476 : < ir !== 'b0000 >");	// Vector No: 869
verify(op === 'b01000000, "Assert 3477 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 3478 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3479 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000100000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 871
#2;

verify(ir === 'b0000, "Assert 3480 : < ir !== 'b0000 >");	// Vector No: 870
verify(op === 'b10000000, "Assert 3481 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3482 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3483 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000100000000000000000000000000:1:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 872
#2;

verify(ir === 'b0000, "Assert 3484 : < ir !== 'b0000 >");	// Vector No: 871
verify(op === 'b00000100, "Assert 3485 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 3486 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3487 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000001000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 873
#2;

verify(ir === 'b0000, "Assert 3488 : < ir !== 'b0000 >");	// Vector No: 872
verify(op === 'b00001000, "Assert 3489 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3490 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3491 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000001000000000000000000000000000:0:1:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 874
#2;

verify(ir === 'b0000, "Assert 3492 : < ir !== 'b0000 >");	// Vector No: 873
verify(op === 'b10000000, "Assert 3493 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3494 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3495 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000001000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 875
#2;

verify(ir === 'b0000, "Assert 3496 : < ir !== 'b0000 >");	// Vector No: 874
verify(op === 'b10000000, "Assert 3497 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3498 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3499 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000001000000000000000000000000000:1:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 876
#2;

verify(ir === 'b0000, "Assert 3500 : < ir !== 'b0000 >");	// Vector No: 875
verify(op === 'b00001000, "Assert 3501 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3502 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3503 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000010000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 877
#2;

verify(ir === 'b0000, "Assert 3504 : < ir !== 'b0000 >");	// Vector No: 876
verify(op === 'b00001000, "Assert 3505 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3506 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3507 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000010000000000000000000000000000:0:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 878
#2;

verify(ir === 'b0001, "Assert 3508 : < ir !== 'b0001 >");	// Vector No: 877
verify(op === 'b00000000, "Assert 3509 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3510 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3511 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000010000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 879
#2;

verify(ir === 'b0000, "Assert 3512 : < ir !== 'b0000 >");	// Vector No: 878
verify(op === 'b10000000, "Assert 3513 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3514 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3515 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000010000000000000000000000000000:1:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 880
#2;

verify(ir === 'b0000, "Assert 3516 : < ir !== 'b0000 >");	// Vector No: 879
verify(op === 'b00010000, "Assert 3517 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 3518 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3519 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000100000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 881
#2;

verify(ir === 'b0000, "Assert 3520 : < ir !== 'b0000 >");	// Vector No: 880
verify(op === 'b00001000, "Assert 3521 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3522 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3523 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000100000000000000000000000000000:0:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 882
#2;

verify(ir === 'b0010, "Assert 3524 : < ir !== 'b0010 >");	// Vector No: 881
verify(op === 'b00000000, "Assert 3525 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3526 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3527 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000100000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 883
#2;

verify(ir === 'b0000, "Assert 3528 : < ir !== 'b0000 >");	// Vector No: 882
verify(op === 'b10000000, "Assert 3529 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3530 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3531 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000100000000000000000000000000000:1:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 884
#2;

verify(ir === 'b0000, "Assert 3532 : < ir !== 'b0000 >");	// Vector No: 883
verify(op === 'b00100000, "Assert 3533 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 3534 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3535 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000001000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 885
#2;

verify(ir === 'b0000, "Assert 3536 : < ir !== 'b0000 >");	// Vector No: 884
verify(op === 'b00001000, "Assert 3537 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3538 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3539 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000001000000000000000000000000000000:0:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 886
#2;

verify(ir === 'b0100, "Assert 3540 : < ir !== 'b0100 >");	// Vector No: 885
verify(op === 'b00000000, "Assert 3541 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3542 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3543 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000001000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 887
#2;

verify(ir === 'b0000, "Assert 3544 : < ir !== 'b0000 >");	// Vector No: 886
verify(op === 'b10000000, "Assert 3545 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3546 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3547 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000001000000000000000000000000000000:1:1:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 888
#2;

verify(ir === 'b0000, "Assert 3548 : < ir !== 'b0000 >");	// Vector No: 887
verify(op === 'b01000000, "Assert 3549 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 3550 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 3551 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000100000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000010000000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 889
#2;

verify(ir === 'b0000, "Assert 3552 : < ir !== 'b0000 >");	// Vector No: 888
verify(op === 'b00001000, "Assert 3553 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3554 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 3555 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000010000000000000000000000100000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 890
#2;

verify(ir === 'b0000, "Assert 3556 : < ir !== 'b0000 >");	// Vector No: 889
verify(op === 'b00000000, "Assert 3557 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3558 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3559 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000100000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 891
#2;

verify(ir === 'b0000, "Assert 3560 : < ir !== 'b0000 >");	// Vector No: 890
verify(op === 'b10000000, "Assert 3561 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3562 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3563 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000100000000000000000000000000000000:1:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 892
#2;

verify(ir === 'b0001, "Assert 3564 : < ir !== 'b0001 >");	// Vector No: 891
verify(op === 'b00000000, "Assert 3565 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3566 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3567 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000001000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000010000000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 893
#2;

verify(ir === 'b0000, "Assert 3568 : < ir !== 'b0000 >");	// Vector No: 892
verify(op === 'b00001000, "Assert 3569 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3570 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 3571 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000010000000000000000000001000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 894
#2;

verify(ir === 'b0000, "Assert 3572 : < ir !== 'b0000 >");	// Vector No: 893
verify(op === 'b00000000, "Assert 3573 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3574 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3575 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000001000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 895
#2;

verify(ir === 'b0000, "Assert 3576 : < ir !== 'b0000 >");	// Vector No: 894
verify(op === 'b10000000, "Assert 3577 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3578 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3579 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000001000000000000000000000000000000000:1:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 896
#2;

verify(ir === 'b0010, "Assert 3580 : < ir !== 'b0010 >");	// Vector No: 895
verify(op === 'b00000000, "Assert 3581 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3582 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3583 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000010000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000010000000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 897
#2;

verify(ir === 'b0000, "Assert 3584 : < ir !== 'b0000 >");	// Vector No: 896
verify(op === 'b00001000, "Assert 3585 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3586 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 3587 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000010000000000000000000010000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 898
#2;

verify(ir === 'b0000, "Assert 3588 : < ir !== 'b0000 >");	// Vector No: 897
verify(op === 'b00000000, "Assert 3589 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3590 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3591 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000010000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 899
#2;

verify(ir === 'b0000, "Assert 3592 : < ir !== 'b0000 >");	// Vector No: 898
verify(op === 'b10000000, "Assert 3593 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3594 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3595 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000010000000000000000000000000000000000:1:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 900
#2;

verify(ir === 'b0100, "Assert 3596 : < ir !== 'b0100 >");	// Vector No: 899
verify(op === 'b00000000, "Assert 3597 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3598 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3599 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000100000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000010000000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 901
#2;

verify(ir === 'b0000, "Assert 3600 : < ir !== 'b0000 >");	// Vector No: 900
verify(op === 'b00001000, "Assert 3601 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3602 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 3603 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000010000000000000000000100000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 902
#2;

verify(ir === 'b0000, "Assert 3604 : < ir !== 'b0000 >");	// Vector No: 901
verify(op === 'b00000000, "Assert 3605 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3606 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3607 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000100000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 903
#2;

verify(ir === 'b0000, "Assert 3608 : < ir !== 'b0000 >");	// Vector No: 902
verify(op === 'b10000000, "Assert 3609 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3610 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3611 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000100000000000000000000000000000000000:1:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 904
#2;

verify(ir === 'b1000, "Assert 3612 : < ir !== 'b1000 >");	// Vector No: 903
verify(op === 'b00000000, "Assert 3613 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3614 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3615 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000001000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000010000000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 905
#2;

verify(ir === 'b0000, "Assert 3616 : < ir !== 'b0000 >");	// Vector No: 904
verify(op === 'b00001000, "Assert 3617 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3618 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 3619 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000010000000000000000001000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 906
#2;

verify(ir === 'b0000, "Assert 3620 : < ir !== 'b0000 >");	// Vector No: 905
verify(op === 'b00000000, "Assert 3621 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3622 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3623 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000001000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000010000000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 907
#2;

verify(ir === 'b0000, "Assert 3624 : < ir !== 'b0000 >");	// Vector No: 906
verify(op === 'b10000000, "Assert 3625 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3626 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 3627 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000010000000000000000001000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 908
#2;

verify(ir === 'b0000, "Assert 3628 : < ir !== 'b0000 >");	// Vector No: 907
verify(op === 'b00000000, "Assert 3629 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3630 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3631 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000010000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000010000000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 909
#2;

verify(ir === 'b0000, "Assert 3632 : < ir !== 'b0000 >");	// Vector No: 908
verify(op === 'b00001000, "Assert 3633 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3634 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 3635 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000010000000000000000010000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 910
#2;

verify(ir === 'b0000, "Assert 3636 : < ir !== 'b0000 >");	// Vector No: 909
verify(op === 'b00000000, "Assert 3637 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3638 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3639 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000010000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000010000000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 911
#2;

verify(ir === 'b0000, "Assert 3640 : < ir !== 'b0000 >");	// Vector No: 910
verify(op === 'b10000000, "Assert 3641 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3642 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 3643 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000010000000000000000010000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 912
#2;

verify(ir === 'b0000, "Assert 3644 : < ir !== 'b0000 >");	// Vector No: 911
verify(op === 'b00000000, "Assert 3645 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3646 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3647 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000100000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000010000000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 913
#2;

verify(ir === 'b0000, "Assert 3648 : < ir !== 'b0000 >");	// Vector No: 912
verify(op === 'b00001000, "Assert 3649 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3650 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 3651 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000010000000000000000100000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 914
#2;

verify(ir === 'b0000, "Assert 3652 : < ir !== 'b0000 >");	// Vector No: 913
verify(op === 'b00000000, "Assert 3653 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3654 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3655 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000100000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000010000000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 915
#2;

verify(ir === 'b0000, "Assert 3656 : < ir !== 'b0000 >");	// Vector No: 914
verify(op === 'b10000000, "Assert 3657 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3658 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 3659 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000010000000000000000100000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 916
#2;

verify(ir === 'b0000, "Assert 3660 : < ir !== 'b0000 >");	// Vector No: 915
verify(op === 'b00000000, "Assert 3661 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3662 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3663 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000001000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000010000000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 917
#2;

verify(ir === 'b0000, "Assert 3664 : < ir !== 'b0000 >");	// Vector No: 916
verify(op === 'b00001000, "Assert 3665 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3666 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 3667 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000010000000000000001000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 918
#2;

verify(ir === 'b0000, "Assert 3668 : < ir !== 'b0000 >");	// Vector No: 917
verify(op === 'b00000000, "Assert 3669 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3670 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3671 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000001000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000010000000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 919
#2;

verify(ir === 'b0000, "Assert 3672 : < ir !== 'b0000 >");	// Vector No: 918
verify(op === 'b10000000, "Assert 3673 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3674 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 3675 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000010000000000000001000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 920
#2;

verify(ir === 'b0000, "Assert 3676 : < ir !== 'b0000 >");	// Vector No: 919
verify(op === 'b00000000, "Assert 3677 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3678 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3679 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000010000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000010000000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 921
#2;

verify(ir === 'b0000, "Assert 3680 : < ir !== 'b0000 >");	// Vector No: 920
verify(op === 'b00001000, "Assert 3681 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3682 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 3683 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000010000000000000010000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 922
#2;

verify(ir === 'b0000, "Assert 3684 : < ir !== 'b0000 >");	// Vector No: 921
verify(op === 'b00000000, "Assert 3685 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3686 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3687 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000010000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000010000000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 923
#2;

verify(ir === 'b0000, "Assert 3688 : < ir !== 'b0000 >");	// Vector No: 922
verify(op === 'b10000000, "Assert 3689 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3690 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 3691 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000010000000000000010000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 924
#2;

verify(ir === 'b0000, "Assert 3692 : < ir !== 'b0000 >");	// Vector No: 923
verify(op === 'b00000000, "Assert 3693 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3694 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3695 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000100000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000010000000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 925
#2;

verify(ir === 'b0000, "Assert 3696 : < ir !== 'b0000 >");	// Vector No: 924
verify(op === 'b00001000, "Assert 3697 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3698 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 3699 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000010000000000000100000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 926
#2;

verify(ir === 'b0000, "Assert 3700 : < ir !== 'b0000 >");	// Vector No: 925
verify(op === 'b00000000, "Assert 3701 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3702 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3703 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000100000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000010000000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 927
#2;

verify(ir === 'b0000, "Assert 3704 : < ir !== 'b0000 >");	// Vector No: 926
verify(op === 'b10000000, "Assert 3705 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3706 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 3707 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000010000000000000100000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 928
#2;

verify(ir === 'b0000, "Assert 3708 : < ir !== 'b0000 >");	// Vector No: 927
verify(op === 'b00000000, "Assert 3709 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3710 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3711 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000001000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000010000000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 929
#2;

verify(ir === 'b0000, "Assert 3712 : < ir !== 'b0000 >");	// Vector No: 928
verify(op === 'b00001000, "Assert 3713 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3714 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 3715 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000010000000000001000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 930
#2;

verify(ir === 'b0000, "Assert 3716 : < ir !== 'b0000 >");	// Vector No: 929
verify(op === 'b00000000, "Assert 3717 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3718 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3719 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000001000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000010000000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 931
#2;

verify(ir === 'b0000, "Assert 3720 : < ir !== 'b0000 >");	// Vector No: 930
verify(op === 'b10000000, "Assert 3721 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3722 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 3723 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000010000000000001000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 932
#2;

verify(ir === 'b0000, "Assert 3724 : < ir !== 'b0000 >");	// Vector No: 931
verify(op === 'b00000000, "Assert 3725 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3726 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3727 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000010000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000010000000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 933
#2;

verify(ir === 'b0000, "Assert 3728 : < ir !== 'b0000 >");	// Vector No: 932
verify(op === 'b00001000, "Assert 3729 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3730 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 3731 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000010000000000010000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 934
#2;

verify(ir === 'b0000, "Assert 3732 : < ir !== 'b0000 >");	// Vector No: 933
verify(op === 'b00000000, "Assert 3733 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3734 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3735 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000010000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000010000000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 935
#2;

verify(ir === 'b0000, "Assert 3736 : < ir !== 'b0000 >");	// Vector No: 934
verify(op === 'b10000000, "Assert 3737 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3738 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 3739 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000010000000000010000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 936
#2;

verify(ir === 'b0000, "Assert 3740 : < ir !== 'b0000 >");	// Vector No: 935
verify(op === 'b00000000, "Assert 3741 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3742 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3743 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000100000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000010000000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 937
#2;

verify(ir === 'b0000, "Assert 3744 : < ir !== 'b0000 >");	// Vector No: 936
verify(op === 'b00001000, "Assert 3745 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3746 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 3747 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000010000000000100000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 938
#2;

verify(ir === 'b0000, "Assert 3748 : < ir !== 'b0000 >");	// Vector No: 937
verify(op === 'b00000000, "Assert 3749 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3750 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3751 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000100000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000010000000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 939
#2;

verify(ir === 'b0000, "Assert 3752 : < ir !== 'b0000 >");	// Vector No: 938
verify(op === 'b10000000, "Assert 3753 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3754 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 3755 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000010000000000100000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 940
#2;

verify(ir === 'b0000, "Assert 3756 : < ir !== 'b0000 >");	// Vector No: 939
verify(op === 'b00000000, "Assert 3757 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3758 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3759 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000001000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000010000000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 941
#2;

verify(ir === 'b0000, "Assert 3760 : < ir !== 'b0000 >");	// Vector No: 940
verify(op === 'b00001000, "Assert 3761 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3762 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 3763 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000010000000001000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 942
#2;

verify(ir === 'b0000, "Assert 3764 : < ir !== 'b0000 >");	// Vector No: 941
verify(op === 'b00000000, "Assert 3765 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3766 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3767 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000001000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000010000000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 943
#2;

verify(ir === 'b0000, "Assert 3768 : < ir !== 'b0000 >");	// Vector No: 942
verify(op === 'b10000000, "Assert 3769 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3770 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 3771 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000010000000001000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 944
#2;

verify(ir === 'b0000, "Assert 3772 : < ir !== 'b0000 >");	// Vector No: 943
verify(op === 'b00000000, "Assert 3773 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3774 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3775 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000010000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000010000000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 945
#2;

verify(ir === 'b0000, "Assert 3776 : < ir !== 'b0000 >");	// Vector No: 944
verify(op === 'b00001000, "Assert 3777 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3778 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 3779 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000010000000010000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 946
#2;

verify(ir === 'b0000, "Assert 3780 : < ir !== 'b0000 >");	// Vector No: 945
verify(op === 'b00000000, "Assert 3781 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3782 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3783 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000010000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000010000000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 947
#2;

verify(ir === 'b0000, "Assert 3784 : < ir !== 'b0000 >");	// Vector No: 946
verify(op === 'b10000000, "Assert 3785 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3786 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 3787 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000010000000010000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 948
#2;

verify(ir === 'b0000, "Assert 3788 : < ir !== 'b0000 >");	// Vector No: 947
verify(op === 'b00000000, "Assert 3789 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3790 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3791 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000100000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000010000000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 949
#2;

verify(ir === 'b0000, "Assert 3792 : < ir !== 'b0000 >");	// Vector No: 948
verify(op === 'b00001000, "Assert 3793 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3794 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 3795 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000010000000100000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 950
#2;

verify(ir === 'b0000, "Assert 3796 : < ir !== 'b0000 >");	// Vector No: 949
verify(op === 'b00000000, "Assert 3797 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3798 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3799 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000100000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000010000000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 951
#2;

verify(ir === 'b0000, "Assert 3800 : < ir !== 'b0000 >");	// Vector No: 950
verify(op === 'b10000000, "Assert 3801 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3802 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 3803 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000010000000100000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 952
#2;

verify(ir === 'b0000, "Assert 3804 : < ir !== 'b0000 >");	// Vector No: 951
verify(op === 'b00000000, "Assert 3805 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3806 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3807 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000001000000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000010000001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 953
#2;

verify(ir === 'b0000, "Assert 3808 : < ir !== 'b0000 >");	// Vector No: 952
verify(op === 'b00001000, "Assert 3809 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3810 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 3811 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000010000001000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 954
#2;

verify(ir === 'b0000, "Assert 3812 : < ir !== 'b0000 >");	// Vector No: 953
verify(op === 'b00000000, "Assert 3813 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3814 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3815 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000001000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000010000001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 955
#2;

verify(ir === 'b0000, "Assert 3816 : < ir !== 'b0000 >");	// Vector No: 954
verify(op === 'b10000000, "Assert 3817 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3818 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 3819 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000010000001000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 956
#2;

verify(ir === 'b0000, "Assert 3820 : < ir !== 'b0000 >");	// Vector No: 955
verify(op === 'b00000000, "Assert 3821 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3822 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3823 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000010000000000000000000000000000000000000000000000000:0:0:0000:00001000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000010000010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 957
#2;

verify(ir === 'b0000, "Assert 3824 : < ir !== 'b0000 >");	// Vector No: 956
verify(op === 'b00001000, "Assert 3825 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3826 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 3827 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000010000010000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 958
#2;

verify(ir === 'b0000, "Assert 3828 : < ir !== 'b0000 >");	// Vector No: 957
verify(op === 'b00000000, "Assert 3829 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3830 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3831 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000010000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000010000010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 959
#2;

verify(ir === 'b0000, "Assert 3832 : < ir !== 'b0000 >");	// Vector No: 958
verify(op === 'b10000000, "Assert 3833 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3834 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 3835 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000010000010000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 960
#2;

verify(ir === 'b0000, "Assert 3836 : < ir !== 'b0000 >");	// Vector No: 959
verify(op === 'b00000000, "Assert 3837 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3838 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3839 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000100000000000000000000000000000000000000000000000000:0:0:0000:00001000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000010000100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 961
#2;

verify(ir === 'b0000, "Assert 3840 : < ir !== 'b0000 >");	// Vector No: 960
verify(op === 'b00001000, "Assert 3841 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3842 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 3843 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000010000100000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 962
#2;

verify(ir === 'b0000, "Assert 3844 : < ir !== 'b0000 >");	// Vector No: 961
verify(op === 'b00000000, "Assert 3845 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3846 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3847 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000100000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000010000100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 963
#2;

verify(ir === 'b0000, "Assert 3848 : < ir !== 'b0000 >");	// Vector No: 962
verify(op === 'b10000000, "Assert 3849 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3850 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 3851 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000010000100000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 964
#2;

verify(ir === 'b0000, "Assert 3852 : < ir !== 'b0000 >");	// Vector No: 963
verify(op === 'b00000000, "Assert 3853 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3854 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3855 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010001000000000000000000000000000000000000000000000000000:0:0:0000:00001000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000010001000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 965
#2;

verify(ir === 'b0000, "Assert 3856 : < ir !== 'b0000 >");	// Vector No: 964
verify(op === 'b00001000, "Assert 3857 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3858 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 3859 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000010001000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010001000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 966
#2;

verify(ir === 'b0000, "Assert 3860 : < ir !== 'b0000 >");	// Vector No: 965
verify(op === 'b00000000, "Assert 3861 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3862 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3863 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010001000000000000000000000000000000000000000000000000000:1:0:0000:10001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010001000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 967
#2;

verify(ir === 'b0000, "Assert 3864 : < ir !== 'b0000 >");	// Vector No: 966
verify(op === 'b10001000, "Assert 3865 : < op !== 'b10001000 >");
verify(extop === 0, "Assert 3866 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3867 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010001000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010001000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 968
#2;

verify(ir === 'b0000, "Assert 3868 : < ir !== 'b0000 >");	// Vector No: 967
verify(op === 'b00000000, "Assert 3869 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3870 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3871 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010010000000000000000000000000000000000000000000000000000:0:0:0000:00001001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010010000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 969
#2;

verify(ir === 'b0000, "Assert 3872 : < ir !== 'b0000 >");	// Vector No: 968
verify(op === 'b00001001, "Assert 3873 : < op !== 'b00001001 >");
verify(extop === 0, "Assert 3874 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3875 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010010000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010010000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 970
#2;

verify(ir === 'b0000, "Assert 3876 : < ir !== 'b0000 >");	// Vector No: 969
verify(op === 'b00000000, "Assert 3877 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3878 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3879 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010010000000000000000000000000000000000000000000000000000:1:0:0000:10010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010010000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 971
#2;

verify(ir === 'b0000, "Assert 3880 : < ir !== 'b0000 >");	// Vector No: 970
verify(op === 'b10010000, "Assert 3881 : < op !== 'b10010000 >");
verify(extop === 0, "Assert 3882 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3883 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010010000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010010000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 972
#2;

verify(ir === 'b0000, "Assert 3884 : < ir !== 'b0000 >");	// Vector No: 971
verify(op === 'b00000000, "Assert 3885 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3886 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3887 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010100000000000000000000000000000000000000000000000000000:0:0:0000:00001010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010100000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 973
#2;

verify(ir === 'b0000, "Assert 3888 : < ir !== 'b0000 >");	// Vector No: 972
verify(op === 'b00001010, "Assert 3889 : < op !== 'b00001010 >");
verify(extop === 0, "Assert 3890 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3891 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010100000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010100000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 974
#2;

verify(ir === 'b0000, "Assert 3892 : < ir !== 'b0000 >");	// Vector No: 973
verify(op === 'b00000000, "Assert 3893 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3894 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3895 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010100000000000000000000000000000000000000000000000000000:1:0:0000:10100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010100000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 975
#2;

verify(ir === 'b0000, "Assert 3896 : < ir !== 'b0000 >");	// Vector No: 974
verify(op === 'b10100000, "Assert 3897 : < op !== 'b10100000 >");
verify(extop === 0, "Assert 3898 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3899 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010100000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010100000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 976
#2;

verify(ir === 'b0000, "Assert 3900 : < ir !== 'b0000 >");	// Vector No: 975
verify(op === 'b00000000, "Assert 3901 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3902 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3903 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000011000000000000000000000000000000000000000000000000000000:0:0:0000:00001100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000011000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 977
#2;

verify(ir === 'b0000, "Assert 3904 : < ir !== 'b0000 >");	// Vector No: 976
verify(op === 'b00001100, "Assert 3905 : < op !== 'b00001100 >");
verify(extop === 0, "Assert 3906 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3907 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000011000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000011000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 978
#2;

verify(ir === 'b0000, "Assert 3908 : < ir !== 'b0000 >");	// Vector No: 977
verify(op === 'b00000000, "Assert 3909 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3910 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3911 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000011000000000000000000000000000000000000000000000000000000:1:0:0000:11000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000011000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 979
#2;

verify(ir === 'b0000, "Assert 3912 : < ir !== 'b0000 >");	// Vector No: 978
verify(op === 'b11000000, "Assert 3913 : < op !== 'b11000000 >");
verify(extop === 0, "Assert 3914 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3915 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000011000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000011000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 980
#2;

verify(ir === 'b0000, "Assert 3916 : < ir !== 'b0000 >");	// Vector No: 979
verify(op === 'b00000000, "Assert 3917 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3918 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3919 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000110000000000000000000000000000000000000000000000000000000:0:0:0000:00011000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000110000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 981
#2;

verify(ir === 'b0000, "Assert 3920 : < ir !== 'b0000 >");	// Vector No: 980
verify(op === 'b00011000, "Assert 3921 : < op !== 'b00011000 >");
verify(extop === 0, "Assert 3922 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3923 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000110000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000110000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 982
#2;

verify(ir === 'b0000, "Assert 3924 : < ir !== 'b0000 >");	// Vector No: 981
verify(op === 'b00000000, "Assert 3925 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3926 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3927 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000110000000000000000000000000000000000000000000000000000000:1:0:0001:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000110000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 983
#2;

verify(ir === 'b0001, "Assert 3928 : < ir !== 'b0001 >");	// Vector No: 982
verify(op === 'b10000000, "Assert 3929 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3930 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3931 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000110000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000110000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 984
#2;

verify(ir === 'b0000, "Assert 3932 : < ir !== 'b0000 >");	// Vector No: 983
verify(op === 'b00000000, "Assert 3933 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3934 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3935 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001010000000000000000000000000000000000000000000000000000000:0:0:0000:00101000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 985
#2;

verify(ir === 'b0000, "Assert 3936 : < ir !== 'b0000 >");	// Vector No: 984
verify(op === 'b00101000, "Assert 3937 : < op !== 'b00101000 >");
verify(extop === 0, "Assert 3938 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3939 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 986
#2;

verify(ir === 'b0000, "Assert 3940 : < ir !== 'b0000 >");	// Vector No: 985
verify(op === 'b00000000, "Assert 3941 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3942 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3943 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001010000000000000000000000000000000000000000000000000000000:1:0:0010:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 987
#2;

verify(ir === 'b0010, "Assert 3944 : < ir !== 'b0010 >");	// Vector No: 986
verify(op === 'b10000000, "Assert 3945 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3946 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3947 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 988
#2;

verify(ir === 'b0000, "Assert 3948 : < ir !== 'b0000 >");	// Vector No: 987
verify(op === 'b00000000, "Assert 3949 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3950 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3951 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010010000000000000000000000000000000000000000000000000000000:0:0:0000:01001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 989
#2;

verify(ir === 'b0000, "Assert 3952 : < ir !== 'b0000 >");	// Vector No: 988
verify(op === 'b01001000, "Assert 3953 : < op !== 'b01001000 >");
verify(extop === 0, "Assert 3954 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3955 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 990
#2;

verify(ir === 'b0000, "Assert 3956 : < ir !== 'b0000 >");	// Vector No: 989
verify(op === 'b00000000, "Assert 3957 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3958 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3959 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010010000000000000000000000000000000000000000000000000000000:1:0:0100:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 991
#2;

verify(ir === 'b0100, "Assert 3960 : < ir !== 'b0100 >");	// Vector No: 990
verify(op === 'b10000000, "Assert 3961 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3962 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3963 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 992
#2;

verify(ir === 'b0000, "Assert 3964 : < ir !== 'b0000 >");	// Vector No: 991
verify(op === 'b00000000, "Assert 3965 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3966 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3967 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100010000000000000000000000000000000000000000000000000000000:0:0:0000:10001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 993
#2;

verify(ir === 'b0000, "Assert 3968 : < ir !== 'b0000 >");	// Vector No: 992
verify(op === 'b10001000, "Assert 3969 : < op !== 'b10001000 >");
verify(extop === 0, "Assert 3970 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3971 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 994
#2;

verify(ir === 'b0000, "Assert 3972 : < ir !== 'b0000 >");	// Vector No: 993
verify(op === 'b00000000, "Assert 3973 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3974 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3975 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100010000000000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 995
#2;

verify(ir === 'b0000, "Assert 3976 : < ir !== 'b0000 >");	// Vector No: 994
verify(op === 'b10000000, "Assert 3977 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3978 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3979 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 996
#2;

verify(ir === 'b0000, "Assert 3980 : < ir !== 'b0000 >");	// Vector No: 995
verify(op === 'b00000000, "Assert 3981 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3982 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3983 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000010000000000000000000000000000000000000000000000000000000:0:0:0001:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 997
#2;

verify(ir === 'b0001, "Assert 3984 : < ir !== 'b0001 >");	// Vector No: 996
verify(op === 'b00001000, "Assert 3985 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 3986 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3987 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 998
#2;

verify(ir === 'b0000, "Assert 3988 : < ir !== 'b0000 >");	// Vector No: 997
verify(op === 'b00000000, "Assert 3989 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3990 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3991 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000010000000000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 999
#2;

verify(ir === 'b0000, "Assert 3992 : < ir !== 'b0000 >");	// Vector No: 998
verify(op === 'b10000000, "Assert 3993 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 3994 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3995 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1000
#2;

verify(ir === 'b0000, "Assert 3996 : < ir !== 'b0000 >");	// Vector No: 999
verify(op === 'b00000000, "Assert 3997 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 3998 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 3999 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000010000000000000000000000000000000000000000000000000000000:0:0:0010:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1001
#2;

verify(ir === 'b0010, "Assert 4000 : < ir !== 'b0010 >");	// Vector No: 1000
verify(op === 'b00001000, "Assert 4001 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 4002 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4003 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1002
#2;

verify(ir === 'b0000, "Assert 4004 : < ir !== 'b0000 >");	// Vector No: 1001
verify(op === 'b00000000, "Assert 4005 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4006 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4007 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000010000000000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1003
#2;

verify(ir === 'b0000, "Assert 4008 : < ir !== 'b0000 >");	// Vector No: 1002
verify(op === 'b10000000, "Assert 4009 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 4010 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4011 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1004
#2;

verify(ir === 'b0000, "Assert 4012 : < ir !== 'b0000 >");	// Vector No: 1003
verify(op === 'b00000000, "Assert 4013 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4014 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4015 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000010000000000000000000000000000000000000000000000000000000:0:0:0100:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1005
#2;

verify(ir === 'b0100, "Assert 4016 : < ir !== 'b0100 >");	// Vector No: 1004
verify(op === 'b00001000, "Assert 4017 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 4018 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4019 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1006
#2;

verify(ir === 'b0000, "Assert 4020 : < ir !== 'b0000 >");	// Vector No: 1005
verify(op === 'b00000000, "Assert 4021 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4022 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4023 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000010000000000000000000000000000000000000000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1007
#2;

verify(ir === 'b0000, "Assert 4024 : < ir !== 'b0000 >");	// Vector No: 1006
verify(op === 'b10000000, "Assert 4025 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 4026 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4027 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1008
#2;

verify(ir === 'b0000, "Assert 4028 : < ir !== 'b0000 >");	// Vector No: 1007
verify(op === 'b00000000, "Assert 4029 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4030 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4031 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000010000000000000000000000000000000000000000000000000000000:0:0:1000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1009
#2;

verify(ir === 'b1000, "Assert 4032 : < ir !== 'b1000 >");	// Vector No: 1008
verify(op === 'b00001000, "Assert 4033 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 4034 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4035 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000010000000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000010000000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1010
#2;

verify(ir === 'b0000, "Assert 4036 : < ir !== 'b0000 >");	// Vector No: 1009
verify(op === 'b00000000, "Assert 4037 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4038 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4039 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000010000000000000000000000000000000000000000000000000000000:1:0:1000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1011
#2;

verify(ir === 'b1000, "Assert 4040 : < ir !== 'b1000 >");	// Vector No: 1010
verify(op === 'b10000000, "Assert 4041 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 4042 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4043 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000010000000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000010000000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1012
#2;

verify(ir === 'b0000, "Assert 4044 : < ir !== 'b0000 >");	// Vector No: 1011
verify(op === 'b00000000, "Assert 4045 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4046 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4047 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000001:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1013
#2;

verify(ir === 'b0000, "Assert 4048 : < ir !== 'b0000 >");	// Vector No: 1012
verify(op === 'b00000000, "Assert 4049 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4050 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4051 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000001:0:1:0000:00000000:1:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1014
#2;

verify(ir === 'b0000, "Assert 4052 : < ir !== 'b0000 >");	// Vector No: 1013
verify(op === 'b00000000, "Assert 4053 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4054 : < extop !== 1 >");
verify(addr === 'b00000000000000000001, "Assert 4055 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000001:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1015
#2;

verify(ir === 'b0000, "Assert 4056 : < ir !== 'b0000 >");	// Vector No: 1014
verify(op === 'b00000000, "Assert 4057 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4058 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4059 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000001:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1016
#2;

verify(ir === 'b0000, "Assert 4060 : < ir !== 'b0000 >");	// Vector No: 1015
verify(op === 'b00000011, "Assert 4061 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4062 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4063 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000001:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1017
#2;

verify(ir === 'b0000, "Assert 4064 : < ir !== 'b0000 >");	// Vector No: 1016
verify(op === 'b00000000, "Assert 4065 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4066 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4067 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000001:0:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000001;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1018
#2;

verify(ir === 'b0000, "Assert 4068 : < ir !== 'b0000 >");	// Vector No: 1017
verify(op === 'b00000000, "Assert 4069 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4070 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 4071 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000001:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1019
#2;

verify(ir === 'b0011, "Assert 4072 : < ir !== 'b0011 >");	// Vector No: 1018
verify(op === 'b11110000, "Assert 4073 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4074 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4075 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000001:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000001;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1020
#2;

verify(ir === 'b0000, "Assert 4076 : < ir !== 'b0000 >");	// Vector No: 1019
verify(op === 'b00000000, "Assert 4077 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4078 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4079 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000010:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1021
#2;

verify(ir === 'b0000, "Assert 4080 : < ir !== 'b0000 >");	// Vector No: 1020
verify(op === 'b00000000, "Assert 4081 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4082 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4083 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000010:0:1:0000:00000000:1:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1022
#2;

verify(ir === 'b0000, "Assert 4084 : < ir !== 'b0000 >");	// Vector No: 1021
verify(op === 'b00000000, "Assert 4085 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4086 : < extop !== 1 >");
verify(addr === 'b00000000000000000010, "Assert 4087 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000010:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1023
#2;

verify(ir === 'b0000, "Assert 4088 : < ir !== 'b0000 >");	// Vector No: 1022
verify(op === 'b00000000, "Assert 4089 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4090 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4091 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000010:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1024
#2;

verify(ir === 'b0000, "Assert 4092 : < ir !== 'b0000 >");	// Vector No: 1023
verify(op === 'b00000011, "Assert 4093 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4094 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4095 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000010:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1025
#2;

verify(ir === 'b0000, "Assert 4096 : < ir !== 'b0000 >");	// Vector No: 1024
verify(op === 'b00000000, "Assert 4097 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4098 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4099 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000010:0:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000010;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1026
#2;

verify(ir === 'b0000, "Assert 4100 : < ir !== 'b0000 >");	// Vector No: 1025
verify(op === 'b00000000, "Assert 4101 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4102 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 4103 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000010:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1027
#2;

verify(ir === 'b0011, "Assert 4104 : < ir !== 'b0011 >");	// Vector No: 1026
verify(op === 'b11110000, "Assert 4105 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4106 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4107 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000010:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000010;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1028
#2;

verify(ir === 'b0000, "Assert 4108 : < ir !== 'b0000 >");	// Vector No: 1027
verify(op === 'b00000000, "Assert 4109 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4110 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4111 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000100:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1029
#2;

verify(ir === 'b0000, "Assert 4112 : < ir !== 'b0000 >");	// Vector No: 1028
verify(op === 'b00000000, "Assert 4113 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4114 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4115 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000100:0:1:0000:00000000:1:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1030
#2;

verify(ir === 'b0000, "Assert 4116 : < ir !== 'b0000 >");	// Vector No: 1029
verify(op === 'b00000000, "Assert 4117 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4118 : < extop !== 1 >");
verify(addr === 'b00000000000000000100, "Assert 4119 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000100:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1031
#2;

verify(ir === 'b0000, "Assert 4120 : < ir !== 'b0000 >");	// Vector No: 1030
verify(op === 'b00000000, "Assert 4121 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4122 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4123 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000100:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1032
#2;

verify(ir === 'b0000, "Assert 4124 : < ir !== 'b0000 >");	// Vector No: 1031
verify(op === 'b00000011, "Assert 4125 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4126 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4127 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000100:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1033
#2;

verify(ir === 'b0000, "Assert 4128 : < ir !== 'b0000 >");	// Vector No: 1032
verify(op === 'b00000000, "Assert 4129 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4130 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4131 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000100:0:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000100;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1034
#2;

verify(ir === 'b0000, "Assert 4132 : < ir !== 'b0000 >");	// Vector No: 1033
verify(op === 'b00000000, "Assert 4133 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4134 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 4135 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000100:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1035
#2;

verify(ir === 'b0011, "Assert 4136 : < ir !== 'b0011 >");	// Vector No: 1034
verify(op === 'b11110000, "Assert 4137 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4138 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4139 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000100:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000100;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1036
#2;

verify(ir === 'b0000, "Assert 4140 : < ir !== 'b0000 >");	// Vector No: 1035
verify(op === 'b00000000, "Assert 4141 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4142 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4143 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000001000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1037
#2;

verify(ir === 'b0000, "Assert 4144 : < ir !== 'b0000 >");	// Vector No: 1036
verify(op === 'b00000000, "Assert 4145 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4146 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4147 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000001000:0:1:0000:00000000:1:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1038
#2;

verify(ir === 'b0000, "Assert 4148 : < ir !== 'b0000 >");	// Vector No: 1037
verify(op === 'b00000000, "Assert 4149 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4150 : < extop !== 1 >");
verify(addr === 'b00000000000000001000, "Assert 4151 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000001000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1039
#2;

verify(ir === 'b0000, "Assert 4152 : < ir !== 'b0000 >");	// Vector No: 1038
verify(op === 'b00000000, "Assert 4153 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4154 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4155 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000001000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1040
#2;

verify(ir === 'b0000, "Assert 4156 : < ir !== 'b0000 >");	// Vector No: 1039
verify(op === 'b00000011, "Assert 4157 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4158 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4159 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000001000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1041
#2;

verify(ir === 'b0000, "Assert 4160 : < ir !== 'b0000 >");	// Vector No: 1040
verify(op === 'b00000000, "Assert 4161 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4162 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4163 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000001000:0:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000001000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1042
#2;

verify(ir === 'b0000, "Assert 4164 : < ir !== 'b0000 >");	// Vector No: 1041
verify(op === 'b00000000, "Assert 4165 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4166 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 4167 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000001000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1043
#2;

verify(ir === 'b0011, "Assert 4168 : < ir !== 'b0011 >");	// Vector No: 1042
verify(op === 'b11110000, "Assert 4169 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4170 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4171 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000001000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000001000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1044
#2;

verify(ir === 'b0000, "Assert 4172 : < ir !== 'b0000 >");	// Vector No: 1043
verify(op === 'b00000000, "Assert 4173 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4174 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4175 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000010000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1045
#2;

verify(ir === 'b0000, "Assert 4176 : < ir !== 'b0000 >");	// Vector No: 1044
verify(op === 'b00000000, "Assert 4177 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4178 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4179 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000010000:0:1:0000:00000000:1:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1046
#2;

verify(ir === 'b0000, "Assert 4180 : < ir !== 'b0000 >");	// Vector No: 1045
verify(op === 'b00000000, "Assert 4181 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4182 : < extop !== 1 >");
verify(addr === 'b00000000000000010000, "Assert 4183 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000010000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1047
#2;

verify(ir === 'b0000, "Assert 4184 : < ir !== 'b0000 >");	// Vector No: 1046
verify(op === 'b00000000, "Assert 4185 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4186 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4187 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000010000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1048
#2;

verify(ir === 'b0000, "Assert 4188 : < ir !== 'b0000 >");	// Vector No: 1047
verify(op === 'b00000011, "Assert 4189 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4190 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4191 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000010000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1049
#2;

verify(ir === 'b0000, "Assert 4192 : < ir !== 'b0000 >");	// Vector No: 1048
verify(op === 'b00000000, "Assert 4193 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4194 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4195 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000010000:0:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000010000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1050
#2;

verify(ir === 'b0000, "Assert 4196 : < ir !== 'b0000 >");	// Vector No: 1049
verify(op === 'b00000000, "Assert 4197 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4198 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 4199 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000010000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1051
#2;

verify(ir === 'b0011, "Assert 4200 : < ir !== 'b0011 >");	// Vector No: 1050
verify(op === 'b11110000, "Assert 4201 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4202 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4203 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000010000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000010000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1052
#2;

verify(ir === 'b0000, "Assert 4204 : < ir !== 'b0000 >");	// Vector No: 1051
verify(op === 'b00000000, "Assert 4205 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4206 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4207 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000100000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1053
#2;

verify(ir === 'b0000, "Assert 4208 : < ir !== 'b0000 >");	// Vector No: 1052
verify(op === 'b00000000, "Assert 4209 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4210 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4211 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000100000:0:1:0000:00000000:1:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1054
#2;

verify(ir === 'b0000, "Assert 4212 : < ir !== 'b0000 >");	// Vector No: 1053
verify(op === 'b00000000, "Assert 4213 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4214 : < extop !== 1 >");
verify(addr === 'b00000000000000100000, "Assert 4215 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000100000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1055
#2;

verify(ir === 'b0000, "Assert 4216 : < ir !== 'b0000 >");	// Vector No: 1054
verify(op === 'b00000000, "Assert 4217 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4218 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4219 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000100000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1056
#2;

verify(ir === 'b0000, "Assert 4220 : < ir !== 'b0000 >");	// Vector No: 1055
verify(op === 'b00000011, "Assert 4221 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4222 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4223 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000100000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1057
#2;

verify(ir === 'b0000, "Assert 4224 : < ir !== 'b0000 >");	// Vector No: 1056
verify(op === 'b00000000, "Assert 4225 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4226 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4227 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000100000:0:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000100000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1058
#2;

verify(ir === 'b0000, "Assert 4228 : < ir !== 'b0000 >");	// Vector No: 1057
verify(op === 'b00000000, "Assert 4229 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4230 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 4231 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000100000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1059
#2;

verify(ir === 'b0011, "Assert 4232 : < ir !== 'b0011 >");	// Vector No: 1058
verify(op === 'b11110000, "Assert 4233 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4234 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4235 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000100000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000100000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1060
#2;

verify(ir === 'b0000, "Assert 4236 : < ir !== 'b0000 >");	// Vector No: 1059
verify(op === 'b00000000, "Assert 4237 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4238 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4239 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000001000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1061
#2;

verify(ir === 'b0000, "Assert 4240 : < ir !== 'b0000 >");	// Vector No: 1060
verify(op === 'b00000000, "Assert 4241 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4242 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4243 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000001000000:0:1:0000:00000000:1:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1062
#2;

verify(ir === 'b0000, "Assert 4244 : < ir !== 'b0000 >");	// Vector No: 1061
verify(op === 'b00000000, "Assert 4245 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4246 : < extop !== 1 >");
verify(addr === 'b00000000000001000000, "Assert 4247 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000001000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1063
#2;

verify(ir === 'b0000, "Assert 4248 : < ir !== 'b0000 >");	// Vector No: 1062
verify(op === 'b00000000, "Assert 4249 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4250 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4251 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000001000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1064
#2;

verify(ir === 'b0000, "Assert 4252 : < ir !== 'b0000 >");	// Vector No: 1063
verify(op === 'b00000011, "Assert 4253 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4254 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4255 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000001000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1065
#2;

verify(ir === 'b0000, "Assert 4256 : < ir !== 'b0000 >");	// Vector No: 1064
verify(op === 'b00000000, "Assert 4257 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4258 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4259 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000001000000:0:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000001000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1066
#2;

verify(ir === 'b0000, "Assert 4260 : < ir !== 'b0000 >");	// Vector No: 1065
verify(op === 'b00000000, "Assert 4261 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4262 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 4263 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000001000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1067
#2;

verify(ir === 'b0011, "Assert 4264 : < ir !== 'b0011 >");	// Vector No: 1066
verify(op === 'b11110000, "Assert 4265 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4266 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4267 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000001000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000001000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1068
#2;

verify(ir === 'b0000, "Assert 4268 : < ir !== 'b0000 >");	// Vector No: 1067
verify(op === 'b00000000, "Assert 4269 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4270 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4271 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000010000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1069
#2;

verify(ir === 'b0000, "Assert 4272 : < ir !== 'b0000 >");	// Vector No: 1068
verify(op === 'b00000000, "Assert 4273 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4274 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4275 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000010000000:0:1:0000:00000000:1:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1070
#2;

verify(ir === 'b0000, "Assert 4276 : < ir !== 'b0000 >");	// Vector No: 1069
verify(op === 'b00000000, "Assert 4277 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4278 : < extop !== 1 >");
verify(addr === 'b00000000000010000000, "Assert 4279 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000010000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1071
#2;

verify(ir === 'b0000, "Assert 4280 : < ir !== 'b0000 >");	// Vector No: 1070
verify(op === 'b00000000, "Assert 4281 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4282 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4283 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000010000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1072
#2;

verify(ir === 'b0000, "Assert 4284 : < ir !== 'b0000 >");	// Vector No: 1071
verify(op === 'b00000011, "Assert 4285 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4286 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4287 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000010000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1073
#2;

verify(ir === 'b0000, "Assert 4288 : < ir !== 'b0000 >");	// Vector No: 1072
verify(op === 'b00000000, "Assert 4289 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4290 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4291 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000010000000:0:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000010000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1074
#2;

verify(ir === 'b0000, "Assert 4292 : < ir !== 'b0000 >");	// Vector No: 1073
verify(op === 'b00000000, "Assert 4293 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4294 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 4295 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000010000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1075
#2;

verify(ir === 'b0011, "Assert 4296 : < ir !== 'b0011 >");	// Vector No: 1074
verify(op === 'b11110000, "Assert 4297 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4298 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4299 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000010000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000010000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1076
#2;

verify(ir === 'b0000, "Assert 4300 : < ir !== 'b0000 >");	// Vector No: 1075
verify(op === 'b00000000, "Assert 4301 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4302 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4303 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000100000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1077
#2;

verify(ir === 'b0000, "Assert 4304 : < ir !== 'b0000 >");	// Vector No: 1076
verify(op === 'b00000000, "Assert 4305 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4306 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4307 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000100000000:0:1:0000:00000000:1:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1078
#2;

verify(ir === 'b0000, "Assert 4308 : < ir !== 'b0000 >");	// Vector No: 1077
verify(op === 'b00000000, "Assert 4309 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4310 : < extop !== 1 >");
verify(addr === 'b00000000000100000000, "Assert 4311 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000100000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1079
#2;

verify(ir === 'b0000, "Assert 4312 : < ir !== 'b0000 >");	// Vector No: 1078
verify(op === 'b00000000, "Assert 4313 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4314 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4315 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000100000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1080
#2;

verify(ir === 'b0000, "Assert 4316 : < ir !== 'b0000 >");	// Vector No: 1079
verify(op === 'b00000011, "Assert 4317 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4318 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4319 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000100000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1081
#2;

verify(ir === 'b0000, "Assert 4320 : < ir !== 'b0000 >");	// Vector No: 1080
verify(op === 'b00000000, "Assert 4321 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4322 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4323 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000100000000:0:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000100000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1082
#2;

verify(ir === 'b0000, "Assert 4324 : < ir !== 'b0000 >");	// Vector No: 1081
verify(op === 'b00000000, "Assert 4325 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4326 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 4327 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000100000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1083
#2;

verify(ir === 'b0011, "Assert 4328 : < ir !== 'b0011 >");	// Vector No: 1082
verify(op === 'b11110000, "Assert 4329 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4330 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4331 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000100000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000100000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1084
#2;

verify(ir === 'b0000, "Assert 4332 : < ir !== 'b0000 >");	// Vector No: 1083
verify(op === 'b00000000, "Assert 4333 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4334 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4335 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000001000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1085
#2;

verify(ir === 'b0000, "Assert 4336 : < ir !== 'b0000 >");	// Vector No: 1084
verify(op === 'b00000000, "Assert 4337 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4338 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4339 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000001000000000:0:1:0000:00000000:1:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1086
#2;

verify(ir === 'b0000, "Assert 4340 : < ir !== 'b0000 >");	// Vector No: 1085
verify(op === 'b00000000, "Assert 4341 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4342 : < extop !== 1 >");
verify(addr === 'b00000000001000000000, "Assert 4343 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000001000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1087
#2;

verify(ir === 'b0000, "Assert 4344 : < ir !== 'b0000 >");	// Vector No: 1086
verify(op === 'b00000000, "Assert 4345 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4346 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4347 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000001000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1088
#2;

verify(ir === 'b0000, "Assert 4348 : < ir !== 'b0000 >");	// Vector No: 1087
verify(op === 'b00000011, "Assert 4349 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4350 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4351 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000001000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1089
#2;

verify(ir === 'b0000, "Assert 4352 : < ir !== 'b0000 >");	// Vector No: 1088
verify(op === 'b00000000, "Assert 4353 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4354 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4355 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000001000000000:0:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000001000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1090
#2;

verify(ir === 'b0000, "Assert 4356 : < ir !== 'b0000 >");	// Vector No: 1089
verify(op === 'b00000000, "Assert 4357 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4358 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 4359 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000001000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1091
#2;

verify(ir === 'b0011, "Assert 4360 : < ir !== 'b0011 >");	// Vector No: 1090
verify(op === 'b11110000, "Assert 4361 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4362 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4363 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000001000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000001000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1092
#2;

verify(ir === 'b0000, "Assert 4364 : < ir !== 'b0000 >");	// Vector No: 1091
verify(op === 'b00000000, "Assert 4365 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4366 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4367 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000010000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1093
#2;

verify(ir === 'b0000, "Assert 4368 : < ir !== 'b0000 >");	// Vector No: 1092
verify(op === 'b00000000, "Assert 4369 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4370 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4371 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000010000000000:0:1:0000:00000000:1:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1094
#2;

verify(ir === 'b0000, "Assert 4372 : < ir !== 'b0000 >");	// Vector No: 1093
verify(op === 'b00000000, "Assert 4373 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4374 : < extop !== 1 >");
verify(addr === 'b00000000010000000000, "Assert 4375 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000010000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1095
#2;

verify(ir === 'b0000, "Assert 4376 : < ir !== 'b0000 >");	// Vector No: 1094
verify(op === 'b00000000, "Assert 4377 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4378 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4379 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000010000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1096
#2;

verify(ir === 'b0000, "Assert 4380 : < ir !== 'b0000 >");	// Vector No: 1095
verify(op === 'b00000011, "Assert 4381 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4382 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4383 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000010000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1097
#2;

verify(ir === 'b0000, "Assert 4384 : < ir !== 'b0000 >");	// Vector No: 1096
verify(op === 'b00000000, "Assert 4385 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4386 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4387 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000010000000000:0:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000010000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1098
#2;

verify(ir === 'b0000, "Assert 4388 : < ir !== 'b0000 >");	// Vector No: 1097
verify(op === 'b00000000, "Assert 4389 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4390 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 4391 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000010000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1099
#2;

verify(ir === 'b0011, "Assert 4392 : < ir !== 'b0011 >");	// Vector No: 1098
verify(op === 'b11110000, "Assert 4393 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4394 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4395 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000010000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000010000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1100
#2;

verify(ir === 'b0000, "Assert 4396 : < ir !== 'b0000 >");	// Vector No: 1099
verify(op === 'b00000000, "Assert 4397 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4398 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4399 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000100000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1101
#2;

verify(ir === 'b0000, "Assert 4400 : < ir !== 'b0000 >");	// Vector No: 1100
verify(op === 'b00000000, "Assert 4401 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4402 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4403 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000100000000000:0:1:0000:00000000:1:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1102
#2;

verify(ir === 'b0000, "Assert 4404 : < ir !== 'b0000 >");	// Vector No: 1101
verify(op === 'b00000000, "Assert 4405 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4406 : < extop !== 1 >");
verify(addr === 'b00000000100000000000, "Assert 4407 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000100000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1103
#2;

verify(ir === 'b0000, "Assert 4408 : < ir !== 'b0000 >");	// Vector No: 1102
verify(op === 'b00000000, "Assert 4409 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4410 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4411 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000100000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1104
#2;

verify(ir === 'b0000, "Assert 4412 : < ir !== 'b0000 >");	// Vector No: 1103
verify(op === 'b00000011, "Assert 4413 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4414 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4415 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000100000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1105
#2;

verify(ir === 'b0000, "Assert 4416 : < ir !== 'b0000 >");	// Vector No: 1104
verify(op === 'b00000000, "Assert 4417 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4418 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4419 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000100000000000:0:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000100000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1106
#2;

verify(ir === 'b0000, "Assert 4420 : < ir !== 'b0000 >");	// Vector No: 1105
verify(op === 'b00000000, "Assert 4421 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4422 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 4423 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000100000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1107
#2;

verify(ir === 'b0011, "Assert 4424 : < ir !== 'b0011 >");	// Vector No: 1106
verify(op === 'b11110000, "Assert 4425 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4426 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4427 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000100000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000100000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1108
#2;

verify(ir === 'b0000, "Assert 4428 : < ir !== 'b0000 >");	// Vector No: 1107
verify(op === 'b00000000, "Assert 4429 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4430 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4431 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000001000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1109
#2;

verify(ir === 'b0000, "Assert 4432 : < ir !== 'b0000 >");	// Vector No: 1108
verify(op === 'b00000000, "Assert 4433 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4434 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4435 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000001000000000000:0:1:0000:00000001:1:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1110
#2;

verify(ir === 'b0000, "Assert 4436 : < ir !== 'b0000 >");	// Vector No: 1109
verify(op === 'b00000001, "Assert 4437 : < op !== 'b00000001 >");
verify(extop === 1, "Assert 4438 : < extop !== 1 >");
verify(addr === 'b00000001000000000000, "Assert 4439 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000001000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1111
#2;

verify(ir === 'b0000, "Assert 4440 : < ir !== 'b0000 >");	// Vector No: 1110
verify(op === 'b00000000, "Assert 4441 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4442 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4443 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000001000000000000:1:1:0000:00000011:0:00000000111100000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1112
#2;

verify(ir === 'b0000, "Assert 4444 : < ir !== 'b0000 >");	// Vector No: 1111
verify(op === 'b00000011, "Assert 4445 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4446 : < extop !== 0 >");
verify(addr === 'b00000000111100000001, "Assert 4447 : < addr !== 'b00000000111100000001 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000001000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1113
#2;

verify(ir === 'b0000, "Assert 4448 : < ir !== 'b0000 >");	// Vector No: 1112
verify(op === 'b00000000, "Assert 4449 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4450 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4451 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000001000000000000:0:1:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000001000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1114
#2;

verify(ir === 'b0000, "Assert 4452 : < ir !== 'b0000 >");	// Vector No: 1113
verify(op === 'b00000000, "Assert 4453 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4454 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 4455 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000001000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1115
#2;

verify(ir === 'b0011, "Assert 4456 : < ir !== 'b0011 >");	// Vector No: 1114
verify(op === 'b11110000, "Assert 4457 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4458 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4459 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000001000000000000:1:1:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000001000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1116
#2;

verify(ir === 'b0000, "Assert 4460 : < ir !== 'b0000 >");	// Vector No: 1115
verify(op === 'b00000000, "Assert 4461 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4462 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 4463 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000010000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1117
#2;

verify(ir === 'b0000, "Assert 4464 : < ir !== 'b0000 >");	// Vector No: 1116
verify(op === 'b00000000, "Assert 4465 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4466 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4467 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000010000000000000:0:1:0000:00000010:1:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1118
#2;

verify(ir === 'b0000, "Assert 4468 : < ir !== 'b0000 >");	// Vector No: 1117
verify(op === 'b00000010, "Assert 4469 : < op !== 'b00000010 >");
verify(extop === 1, "Assert 4470 : < extop !== 1 >");
verify(addr === 'b00000010000000000000, "Assert 4471 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000010000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1119
#2;

verify(ir === 'b0000, "Assert 4472 : < ir !== 'b0000 >");	// Vector No: 1118
verify(op === 'b00000000, "Assert 4473 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4474 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4475 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000010000000000000:1:1:0000:00000011:0:00000000111100000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1120
#2;

verify(ir === 'b0000, "Assert 4476 : < ir !== 'b0000 >");	// Vector No: 1119
verify(op === 'b00000011, "Assert 4477 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4478 : < extop !== 0 >");
verify(addr === 'b00000000111100000010, "Assert 4479 : < addr !== 'b00000000111100000010 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000010000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1121
#2;

verify(ir === 'b0000, "Assert 4480 : < ir !== 'b0000 >");	// Vector No: 1120
verify(op === 'b00000000, "Assert 4481 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4482 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4483 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000010000000000000:0:1:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000010000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1122
#2;

verify(ir === 'b0000, "Assert 4484 : < ir !== 'b0000 >");	// Vector No: 1121
verify(op === 'b00000000, "Assert 4485 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4486 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 4487 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000010000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1123
#2;

verify(ir === 'b0011, "Assert 4488 : < ir !== 'b0011 >");	// Vector No: 1122
verify(op === 'b11110000, "Assert 4489 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4490 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4491 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000010000000000000:1:1:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000010000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1124
#2;

verify(ir === 'b0000, "Assert 4492 : < ir !== 'b0000 >");	// Vector No: 1123
verify(op === 'b00000000, "Assert 4493 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4494 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 4495 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000100000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1125
#2;

verify(ir === 'b0000, "Assert 4496 : < ir !== 'b0000 >");	// Vector No: 1124
verify(op === 'b00000000, "Assert 4497 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4498 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4499 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000100000000000000:0:1:0000:00000100:1:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1126
#2;

verify(ir === 'b0000, "Assert 4500 : < ir !== 'b0000 >");	// Vector No: 1125
verify(op === 'b00000100, "Assert 4501 : < op !== 'b00000100 >");
verify(extop === 1, "Assert 4502 : < extop !== 1 >");
verify(addr === 'b00000100000000000000, "Assert 4503 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000100000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1127
#2;

verify(ir === 'b0000, "Assert 4504 : < ir !== 'b0000 >");	// Vector No: 1126
verify(op === 'b00000000, "Assert 4505 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4506 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4507 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000100000000000000:1:1:0000:00000011:0:00000000111100000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1128
#2;

verify(ir === 'b0000, "Assert 4508 : < ir !== 'b0000 >");	// Vector No: 1127
verify(op === 'b00000011, "Assert 4509 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4510 : < extop !== 0 >");
verify(addr === 'b00000000111100000100, "Assert 4511 : < addr !== 'b00000000111100000100 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000100000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1129
#2;

verify(ir === 'b0000, "Assert 4512 : < ir !== 'b0000 >");	// Vector No: 1128
verify(op === 'b00000000, "Assert 4513 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4514 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4515 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000100000000000000:0:1:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000100000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1130
#2;

verify(ir === 'b0000, "Assert 4516 : < ir !== 'b0000 >");	// Vector No: 1129
verify(op === 'b00000000, "Assert 4517 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4518 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 4519 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000100000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1131
#2;

verify(ir === 'b0011, "Assert 4520 : < ir !== 'b0011 >");	// Vector No: 1130
verify(op === 'b11110000, "Assert 4521 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4522 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4523 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000100000000000000:1:1:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000100000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1132
#2;

verify(ir === 'b0000, "Assert 4524 : < ir !== 'b0000 >");	// Vector No: 1131
verify(op === 'b00000000, "Assert 4525 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4526 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 4527 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100001000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100001000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1133
#2;

verify(ir === 'b0000, "Assert 4528 : < ir !== 'b0000 >");	// Vector No: 1132
verify(op === 'b00000000, "Assert 4529 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4530 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4531 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100001000000000000000:0:1:0000:00001000:1:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100001000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1134
#2;

verify(ir === 'b0000, "Assert 4532 : < ir !== 'b0000 >");	// Vector No: 1133
verify(op === 'b00001000, "Assert 4533 : < op !== 'b00001000 >");
verify(extop === 1, "Assert 4534 : < extop !== 1 >");
verify(addr === 'b00001000000000000000, "Assert 4535 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100001000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100001000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1135
#2;

verify(ir === 'b0000, "Assert 4536 : < ir !== 'b0000 >");	// Vector No: 1134
verify(op === 'b00000000, "Assert 4537 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4538 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4539 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100001000000000000000:1:1:0000:00000011:0:00000000111100001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100001000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1136
#2;

verify(ir === 'b0000, "Assert 4540 : < ir !== 'b0000 >");	// Vector No: 1135
verify(op === 'b00000011, "Assert 4541 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4542 : < extop !== 0 >");
verify(addr === 'b00000000111100001000, "Assert 4543 : < addr !== 'b00000000111100001000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000001000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1137
#2;

verify(ir === 'b0000, "Assert 4544 : < ir !== 'b0000 >");	// Vector No: 1136
verify(op === 'b00000000, "Assert 4545 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4546 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4547 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000001000000000000000:0:1:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000001000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1138
#2;

verify(ir === 'b0000, "Assert 4548 : < ir !== 'b0000 >");	// Vector No: 1137
verify(op === 'b00000000, "Assert 4549 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4550 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 4551 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000001000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1139
#2;

verify(ir === 'b0011, "Assert 4552 : < ir !== 'b0011 >");	// Vector No: 1138
verify(op === 'b11110000, "Assert 4553 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4554 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4555 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000001000000000000000:1:1:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000001000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1140
#2;

verify(ir === 'b0000, "Assert 4556 : < ir !== 'b0000 >");	// Vector No: 1139
verify(op === 'b00000000, "Assert 4557 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4558 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 4559 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100010000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100010000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1141
#2;

verify(ir === 'b0000, "Assert 4560 : < ir !== 'b0000 >");	// Vector No: 1140
verify(op === 'b00000000, "Assert 4561 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4562 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4563 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100010000000000000000:0:1:0000:00010000:1:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100010000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1142
#2;

verify(ir === 'b0000, "Assert 4564 : < ir !== 'b0000 >");	// Vector No: 1141
verify(op === 'b00010000, "Assert 4565 : < op !== 'b00010000 >");
verify(extop === 1, "Assert 4566 : < extop !== 1 >");
verify(addr === 'b00010000000000000000, "Assert 4567 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100010000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100010000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1143
#2;

verify(ir === 'b0000, "Assert 4568 : < ir !== 'b0000 >");	// Vector No: 1142
verify(op === 'b00000000, "Assert 4569 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4570 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4571 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100010000000000000000:1:1:0000:00000011:0:00000000111100010000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100010000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1144
#2;

verify(ir === 'b0000, "Assert 4572 : < ir !== 'b0000 >");	// Vector No: 1143
verify(op === 'b00000011, "Assert 4573 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4574 : < extop !== 0 >");
verify(addr === 'b00000000111100010000, "Assert 4575 : < addr !== 'b00000000111100010000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000010000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1145
#2;

verify(ir === 'b0000, "Assert 4576 : < ir !== 'b0000 >");	// Vector No: 1144
verify(op === 'b00000000, "Assert 4577 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4578 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4579 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000010000000000000000:0:1:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000010000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1146
#2;

verify(ir === 'b0000, "Assert 4580 : < ir !== 'b0000 >");	// Vector No: 1145
verify(op === 'b00000000, "Assert 4581 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4582 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 4583 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000010000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1147
#2;

verify(ir === 'b0011, "Assert 4584 : < ir !== 'b0011 >");	// Vector No: 1146
verify(op === 'b11110000, "Assert 4585 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4586 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4587 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000010000000000000000:1:1:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000010000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1148
#2;

verify(ir === 'b0000, "Assert 4588 : < ir !== 'b0000 >");	// Vector No: 1147
verify(op === 'b00000000, "Assert 4589 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4590 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 4591 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100100000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100100000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1149
#2;

verify(ir === 'b0000, "Assert 4592 : < ir !== 'b0000 >");	// Vector No: 1148
verify(op === 'b00000000, "Assert 4593 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4594 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4595 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100100000000000000000:0:1:0000:00100000:1:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100100000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1150
#2;

verify(ir === 'b0000, "Assert 4596 : < ir !== 'b0000 >");	// Vector No: 1149
verify(op === 'b00100000, "Assert 4597 : < op !== 'b00100000 >");
verify(extop === 1, "Assert 4598 : < extop !== 1 >");
verify(addr === 'b00100000000000000000, "Assert 4599 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100100000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100100000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1151
#2;

verify(ir === 'b0000, "Assert 4600 : < ir !== 'b0000 >");	// Vector No: 1150
verify(op === 'b00000000, "Assert 4601 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4602 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4603 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100100000000000000000:1:1:0000:00000011:0:00000000111100100000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100100000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1152
#2;

verify(ir === 'b0000, "Assert 4604 : < ir !== 'b0000 >");	// Vector No: 1151
verify(op === 'b00000011, "Assert 4605 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4606 : < extop !== 0 >");
verify(addr === 'b00000000111100100000, "Assert 4607 : < addr !== 'b00000000111100100000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000100000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1153
#2;

verify(ir === 'b0000, "Assert 4608 : < ir !== 'b0000 >");	// Vector No: 1152
verify(op === 'b00000000, "Assert 4609 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4610 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4611 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000100000000000000000:0:1:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000100000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1154
#2;

verify(ir === 'b0000, "Assert 4612 : < ir !== 'b0000 >");	// Vector No: 1153
verify(op === 'b00000000, "Assert 4613 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4614 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 4615 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000100000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1155
#2;

verify(ir === 'b0011, "Assert 4616 : < ir !== 'b0011 >");	// Vector No: 1154
verify(op === 'b11110000, "Assert 4617 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4618 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4619 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000100000000000000000:1:1:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000100000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1156
#2;

verify(ir === 'b0000, "Assert 4620 : < ir !== 'b0000 >");	// Vector No: 1155
verify(op === 'b00000000, "Assert 4621 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4622 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 4623 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111101000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111101000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1157
#2;

verify(ir === 'b0000, "Assert 4624 : < ir !== 'b0000 >");	// Vector No: 1156
verify(op === 'b00000000, "Assert 4625 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4626 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4627 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111101000000000000000000:0:1:0000:01000000:1:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111101000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1158
#2;

verify(ir === 'b0000, "Assert 4628 : < ir !== 'b0000 >");	// Vector No: 1157
verify(op === 'b01000000, "Assert 4629 : < op !== 'b01000000 >");
verify(extop === 1, "Assert 4630 : < extop !== 1 >");
verify(addr === 'b01000000000000000000, "Assert 4631 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111101000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111101000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1159
#2;

verify(ir === 'b0000, "Assert 4632 : < ir !== 'b0000 >");	// Vector No: 1158
verify(op === 'b00000000, "Assert 4633 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4634 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4635 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111101000000000000000000:1:1:0000:00000011:0:00000000111101000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111101000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1160
#2;

verify(ir === 'b0000, "Assert 4636 : < ir !== 'b0000 >");	// Vector No: 1159
verify(op === 'b00000011, "Assert 4637 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4638 : < extop !== 0 >");
verify(addr === 'b00000000111101000000, "Assert 4639 : < addr !== 'b00000000111101000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000001000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1161
#2;

verify(ir === 'b0000, "Assert 4640 : < ir !== 'b0000 >");	// Vector No: 1160
verify(op === 'b00000000, "Assert 4641 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4642 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4643 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000001000000000000000000:0:1:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000001000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1162
#2;

verify(ir === 'b0000, "Assert 4644 : < ir !== 'b0000 >");	// Vector No: 1161
verify(op === 'b00000000, "Assert 4645 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4646 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 4647 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000001000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1163
#2;

verify(ir === 'b0011, "Assert 4648 : < ir !== 'b0011 >");	// Vector No: 1162
verify(op === 'b11110000, "Assert 4649 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4650 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4651 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000001000000000000000000:1:1:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000001000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1164
#2;

verify(ir === 'b0000, "Assert 4652 : < ir !== 'b0000 >");	// Vector No: 1163
verify(op === 'b00000000, "Assert 4653 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4654 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 4655 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111110000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111110000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1165
#2;

verify(ir === 'b0000, "Assert 4656 : < ir !== 'b0000 >");	// Vector No: 1164
verify(op === 'b00000000, "Assert 4657 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4658 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4659 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111110000000000000000000:0:1:0000:10000000:1:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111110000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1166
#2;

verify(ir === 'b0000, "Assert 4660 : < ir !== 'b0000 >");	// Vector No: 1165
verify(op === 'b10000000, "Assert 4661 : < op !== 'b10000000 >");
verify(extop === 1, "Assert 4662 : < extop !== 1 >");
verify(addr === 'b10000000000000000000, "Assert 4663 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111110000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111110000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1167
#2;

verify(ir === 'b0000, "Assert 4664 : < ir !== 'b0000 >");	// Vector No: 1166
verify(op === 'b00000000, "Assert 4665 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4666 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4667 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111110000000000000000000:1:1:0000:00000011:0:00000000111110000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111110000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1168
#2;

verify(ir === 'b0000, "Assert 4668 : < ir !== 'b0000 >");	// Vector No: 1167
verify(op === 'b00000011, "Assert 4669 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4670 : < extop !== 0 >");
verify(addr === 'b00000000111110000000, "Assert 4671 : < addr !== 'b00000000111110000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000010000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1169
#2;

verify(ir === 'b0000, "Assert 4672 : < ir !== 'b0000 >");	// Vector No: 1168
verify(op === 'b00000000, "Assert 4673 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4674 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4675 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000010000000000000000000:0:1:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000010000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1170
#2;

verify(ir === 'b0000, "Assert 4676 : < ir !== 'b0000 >");	// Vector No: 1169
verify(op === 'b00000000, "Assert 4677 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4678 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 4679 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000010000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1171
#2;

verify(ir === 'b0011, "Assert 4680 : < ir !== 'b0011 >");	// Vector No: 1170
verify(op === 'b11110000, "Assert 4681 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4682 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4683 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000010000000000000000000:1:1:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000010000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1172
#2;

verify(ir === 'b0000, "Assert 4684 : < ir !== 'b0000 >");	// Vector No: 1171
verify(op === 'b00000000, "Assert 4685 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4686 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 4687 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1173
#2;

verify(ir === 'b0000, "Assert 4688 : < ir !== 'b0000 >");	// Vector No: 1172
verify(op === 'b00000000, "Assert 4689 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4690 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4691 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1174
#2;

verify(ir === 'b0000, "Assert 4692 : < ir !== 'b0000 >");	// Vector No: 1173
verify(op === 'b00000000, "Assert 4693 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4694 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4695 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1175
#2;

verify(ir === 'b0000, "Assert 4696 : < ir !== 'b0000 >");	// Vector No: 1174
verify(op === 'b00000000, "Assert 4697 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4698 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4699 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1176
#2;

verify(ir === 'b0000, "Assert 4700 : < ir !== 'b0000 >");	// Vector No: 1175
verify(op === 'b00000011, "Assert 4701 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4702 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4703 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000100000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1177
#2;

verify(ir === 'b0000, "Assert 4704 : < ir !== 'b0000 >");	// Vector No: 1176
verify(op === 'b00000000, "Assert 4705 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4706 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4707 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000100000000000000000000:0:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1178
#2;

verify(ir === 'b0000, "Assert 4708 : < ir !== 'b0000 >");	// Vector No: 1177
verify(op === 'b00000001, "Assert 4709 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 4710 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4711 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000100000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1179
#2;

verify(ir === 'b0011, "Assert 4712 : < ir !== 'b0011 >");	// Vector No: 1178
verify(op === 'b11110000, "Assert 4713 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4714 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4715 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000100000000000000000000:1:1:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1180
#2;

verify(ir === 'b0000, "Assert 4716 : < ir !== 'b0000 >");	// Vector No: 1179
verify(op === 'b00000000, "Assert 4717 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4718 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 4719 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000001000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1181
#2;

verify(ir === 'b0000, "Assert 4720 : < ir !== 'b0000 >");	// Vector No: 1180
verify(op === 'b00000000, "Assert 4721 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4722 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4723 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000001000000000000000000000:0:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000001000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1182
#2;

verify(ir === 'b0000, "Assert 4724 : < ir !== 'b0000 >");	// Vector No: 1181
verify(op === 'b00000010, "Assert 4725 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 4726 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4727 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000001000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1183
#2;

verify(ir === 'b0011, "Assert 4728 : < ir !== 'b0011 >");	// Vector No: 1182
verify(op === 'b11110000, "Assert 4729 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4730 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4731 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000001000000000000000000000:1:1:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000001000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1184
#2;

verify(ir === 'b0000, "Assert 4732 : < ir !== 'b0000 >");	// Vector No: 1183
verify(op === 'b00000000, "Assert 4733 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4734 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 4735 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000010000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1185
#2;

verify(ir === 'b0000, "Assert 4736 : < ir !== 'b0000 >");	// Vector No: 1184
verify(op === 'b00000000, "Assert 4737 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4738 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4739 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000010000000000000000000000:0:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000010000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1186
#2;

verify(ir === 'b0000, "Assert 4740 : < ir !== 'b0000 >");	// Vector No: 1185
verify(op === 'b00000100, "Assert 4741 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 4742 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4743 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000010000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1187
#2;

verify(ir === 'b0011, "Assert 4744 : < ir !== 'b0011 >");	// Vector No: 1186
verify(op === 'b11110000, "Assert 4745 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4746 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4747 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000010000000000000000000000:1:1:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000010000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1188
#2;

verify(ir === 'b0000, "Assert 4748 : < ir !== 'b0000 >");	// Vector No: 1187
verify(op === 'b00000000, "Assert 4749 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4750 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 4751 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000100000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1189
#2;

verify(ir === 'b0000, "Assert 4752 : < ir !== 'b0000 >");	// Vector No: 1188
verify(op === 'b00000000, "Assert 4753 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4754 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4755 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000100000000000000000000000:0:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000100000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1190
#2;

verify(ir === 'b0000, "Assert 4756 : < ir !== 'b0000 >");	// Vector No: 1189
verify(op === 'b00001000, "Assert 4757 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 4758 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4759 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000100000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1191
#2;

verify(ir === 'b0011, "Assert 4760 : < ir !== 'b0011 >");	// Vector No: 1190
verify(op === 'b11110000, "Assert 4761 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4762 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4763 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000100000000000000000000000:1:1:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000100000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1192
#2;

verify(ir === 'b0000, "Assert 4764 : < ir !== 'b0000 >");	// Vector No: 1191
verify(op === 'b00000000, "Assert 4765 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4766 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 4767 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000001000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1193
#2;

verify(ir === 'b0000, "Assert 4768 : < ir !== 'b0000 >");	// Vector No: 1192
verify(op === 'b00000000, "Assert 4769 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4770 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4771 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000001000000000000000000000000:0:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000001000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1194
#2;

verify(ir === 'b0000, "Assert 4772 : < ir !== 'b0000 >");	// Vector No: 1193
verify(op === 'b00010000, "Assert 4773 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 4774 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4775 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000001000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1195
#2;

verify(ir === 'b0011, "Assert 4776 : < ir !== 'b0011 >");	// Vector No: 1194
verify(op === 'b11110000, "Assert 4777 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4778 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4779 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000001000000000000000000000000:1:1:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000001000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1196
#2;

verify(ir === 'b0000, "Assert 4780 : < ir !== 'b0000 >");	// Vector No: 1195
verify(op === 'b00000001, "Assert 4781 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 4782 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4783 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000010000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1197
#2;

verify(ir === 'b0000, "Assert 4784 : < ir !== 'b0000 >");	// Vector No: 1196
verify(op === 'b00000000, "Assert 4785 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4786 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4787 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000010000000000000000000000000:0:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000010000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1198
#2;

verify(ir === 'b0000, "Assert 4788 : < ir !== 'b0000 >");	// Vector No: 1197
verify(op === 'b00100000, "Assert 4789 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 4790 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4791 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000010000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1199
#2;

verify(ir === 'b0011, "Assert 4792 : < ir !== 'b0011 >");	// Vector No: 1198
verify(op === 'b11110000, "Assert 4793 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4794 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4795 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000010000000000000000000000000:1:1:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000010000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1200
#2;

verify(ir === 'b0000, "Assert 4796 : < ir !== 'b0000 >");	// Vector No: 1199
verify(op === 'b00000010, "Assert 4797 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 4798 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4799 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000100000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1201
#2;

verify(ir === 'b0000, "Assert 4800 : < ir !== 'b0000 >");	// Vector No: 1200
verify(op === 'b00000000, "Assert 4801 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4802 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4803 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000100000000000000000000000000:0:1:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000100000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1202
#2;

verify(ir === 'b0000, "Assert 4804 : < ir !== 'b0000 >");	// Vector No: 1201
verify(op === 'b01000000, "Assert 4805 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 4806 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4807 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000100000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1203
#2;

verify(ir === 'b0011, "Assert 4808 : < ir !== 'b0011 >");	// Vector No: 1202
verify(op === 'b11110000, "Assert 4809 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4810 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4811 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000100000000000000000000000000:1:1:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000100000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1204
#2;

verify(ir === 'b0000, "Assert 4812 : < ir !== 'b0000 >");	// Vector No: 1203
verify(op === 'b00000100, "Assert 4813 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 4814 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4815 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000001000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1205
#2;

verify(ir === 'b0000, "Assert 4816 : < ir !== 'b0000 >");	// Vector No: 1204
verify(op === 'b00000000, "Assert 4817 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4818 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4819 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000001000000000000000000000000000:0:1:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000001000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1206
#2;

verify(ir === 'b0000, "Assert 4820 : < ir !== 'b0000 >");	// Vector No: 1205
verify(op === 'b10000000, "Assert 4821 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 4822 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4823 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000001000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1207
#2;

verify(ir === 'b0011, "Assert 4824 : < ir !== 'b0011 >");	// Vector No: 1206
verify(op === 'b11110000, "Assert 4825 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4826 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4827 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000001000000000000000000000000000:1:1:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000001000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1208
#2;

verify(ir === 'b0000, "Assert 4828 : < ir !== 'b0000 >");	// Vector No: 1207
verify(op === 'b00001000, "Assert 4829 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 4830 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4831 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010011111100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1209
#2;

verify(ir === 'b0000, "Assert 4832 : < ir !== 'b0000 >");	// Vector No: 1208
verify(op === 'b00000000, "Assert 4833 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4834 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4835 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010011111100000000000000000000:0:1:0001:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1210
#2;

verify(ir === 'b0001, "Assert 4836 : < ir !== 'b0001 >");	// Vector No: 1209
verify(op === 'b00000000, "Assert 4837 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4838 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4839 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1211
#2;

verify(ir === 'b0000, "Assert 4840 : < ir !== 'b0000 >");	// Vector No: 1210
verify(op === 'b00000000, "Assert 4841 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4842 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4843 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000010011111100000000000000000000:1:1:0000:00010011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000010011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1212
#2;

verify(ir === 'b0000, "Assert 4844 : < ir !== 'b0000 >");	// Vector No: 1211
verify(op === 'b00010011, "Assert 4845 : < op !== 'b00010011 >");
verify(extop === 0, "Assert 4846 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4847 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000010000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1213
#2;

verify(ir === 'b0000, "Assert 4848 : < ir !== 'b0000 >");	// Vector No: 1212
verify(op === 'b00000000, "Assert 4849 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4850 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4851 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000010000000000000000000000000000:0:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000010000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1214
#2;

verify(ir === 'b0001, "Assert 4852 : < ir !== 'b0001 >");	// Vector No: 1213
verify(op === 'b00000000, "Assert 4853 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4854 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4855 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000010000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1215
#2;

verify(ir === 'b0011, "Assert 4856 : < ir !== 'b0011 >");	// Vector No: 1214
verify(op === 'b11110000, "Assert 4857 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4858 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4859 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000010000000000000000000000000000:1:1:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000010000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1216
#2;

verify(ir === 'b0000, "Assert 4860 : < ir !== 'b0000 >");	// Vector No: 1215
verify(op === 'b00010000, "Assert 4861 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 4862 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4863 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100011111100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1217
#2;

verify(ir === 'b0000, "Assert 4864 : < ir !== 'b0000 >");	// Vector No: 1216
verify(op === 'b00000000, "Assert 4865 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4866 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4867 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100011111100000000000000000000:0:1:0010:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1218
#2;

verify(ir === 'b0010, "Assert 4868 : < ir !== 'b0010 >");	// Vector No: 1217
verify(op === 'b00000000, "Assert 4869 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4870 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4871 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1219
#2;

verify(ir === 'b0000, "Assert 4872 : < ir !== 'b0000 >");	// Vector No: 1218
verify(op === 'b00000000, "Assert 4873 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4874 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4875 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000000100011111100000000000000000000:1:1:0000:00100011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000000100011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1220
#2;

verify(ir === 'b0000, "Assert 4876 : < ir !== 'b0000 >");	// Vector No: 1219
verify(op === 'b00100011, "Assert 4877 : < op !== 'b00100011 >");
verify(extop === 0, "Assert 4878 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4879 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000100000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1221
#2;

verify(ir === 'b0000, "Assert 4880 : < ir !== 'b0000 >");	// Vector No: 1220
verify(op === 'b00000000, "Assert 4881 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4882 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4883 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000100000000000000000000000000000:0:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000100000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1222
#2;

verify(ir === 'b0010, "Assert 4884 : < ir !== 'b0010 >");	// Vector No: 1221
verify(op === 'b00000000, "Assert 4885 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4886 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4887 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000100000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1223
#2;

verify(ir === 'b0011, "Assert 4888 : < ir !== 'b0011 >");	// Vector No: 1222
verify(op === 'b11110000, "Assert 4889 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4890 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4891 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000100000000000000000000000000000:1:1:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000100000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1224
#2;

verify(ir === 'b0000, "Assert 4892 : < ir !== 'b0000 >");	// Vector No: 1223
verify(op === 'b00100000, "Assert 4893 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 4894 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4895 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1225
#2;

verify(ir === 'b0000, "Assert 4896 : < ir !== 'b0000 >");	// Vector No: 1224
verify(op === 'b00000000, "Assert 4897 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4898 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4899 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000011111100000000000000000000:0:1:0100:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1226
#2;

verify(ir === 'b0100, "Assert 4900 : < ir !== 'b0100 >");	// Vector No: 1225
verify(op === 'b00000000, "Assert 4901 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4902 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4903 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1227
#2;

verify(ir === 'b0000, "Assert 4904 : < ir !== 'b0000 >");	// Vector No: 1226
verify(op === 'b00000000, "Assert 4905 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4906 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4907 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000001000011111100000000000000000000:1:1:0000:01000011:0:00000111111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000001000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1228
#2;

verify(ir === 'b0000, "Assert 4908 : < ir !== 'b0000 >");	// Vector No: 1227
verify(op === 'b01000011, "Assert 4909 : < op !== 'b01000011 >");
verify(extop === 0, "Assert 4910 : < extop !== 0 >");
verify(addr === 'b00000111111100000000, "Assert 4911 : < addr !== 'b00000111111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000001000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1229
#2;

verify(ir === 'b0000, "Assert 4912 : < ir !== 'b0000 >");	// Vector No: 1228
verify(op === 'b00000000, "Assert 4913 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4914 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4915 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000001000000000000000000000000000000:0:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000001000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1230
#2;

verify(ir === 'b0100, "Assert 4916 : < ir !== 'b0100 >");	// Vector No: 1229
verify(op === 'b00000000, "Assert 4917 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4918 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4919 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000001000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1231
#2;

verify(ir === 'b0011, "Assert 4920 : < ir !== 'b0011 >");	// Vector No: 1230
verify(op === 'b11110000, "Assert 4921 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4922 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4923 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000001000000000000000000000000000000:1:1:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000001000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1232
#2;

verify(ir === 'b0000, "Assert 4924 : < ir !== 'b0000 >");	// Vector No: 1231
verify(op === 'b01000000, "Assert 4925 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 4926 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 4927 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1233
#2;

verify(ir === 'b0000, "Assert 4928 : < ir !== 'b0000 >");	// Vector No: 1232
verify(op === 'b00000000, "Assert 4929 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4930 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4931 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000011111100000000000000000000:0:1:1000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1234
#2;

verify(ir === 'b1000, "Assert 4932 : < ir !== 'b1000 >");	// Vector No: 1233
verify(op === 'b00000000, "Assert 4933 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4934 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4935 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1235
#2;

verify(ir === 'b0000, "Assert 4936 : < ir !== 'b0000 >");	// Vector No: 1234
verify(op === 'b00000000, "Assert 4937 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4938 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4939 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000010000011111100000000000000000000:1:1:0000:00000000:0:00000011111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000010000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1236
#2;

verify(ir === 'b0000, "Assert 4940 : < ir !== 'b0000 >");	// Vector No: 1235
verify(op === 'b00000000, "Assert 4941 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4942 : < extop !== 0 >");
verify(addr === 'b00000011111100000000, "Assert 4943 : < addr !== 'b00000011111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000010000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1237
#2;

verify(ir === 'b0000, "Assert 4944 : < ir !== 'b0000 >");	// Vector No: 1236
verify(op === 'b00000000, "Assert 4945 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4946 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4947 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000010000000000000000000000000000000:0:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000010000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1238
#2;

verify(ir === 'b1000, "Assert 4948 : < ir !== 'b1000 >");	// Vector No: 1237
verify(op === 'b00000000, "Assert 4949 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4950 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4951 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000010000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1239
#2;

verify(ir === 'b0011, "Assert 4952 : < ir !== 'b0011 >");	// Vector No: 1238
verify(op === 'b11110000, "Assert 4953 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4954 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4955 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000010000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000010000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1240
#2;

verify(ir === 'b0000, "Assert 4956 : < ir !== 'b0000 >");	// Vector No: 1239
verify(op === 'b00000000, "Assert 4957 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4958 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4959 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1241
#2;

verify(ir === 'b0000, "Assert 4960 : < ir !== 'b0000 >");	// Vector No: 1240
verify(op === 'b00000000, "Assert 4961 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4962 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 4963 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1242
#2;

verify(ir === 'b0000, "Assert 4964 : < ir !== 'b0000 >");	// Vector No: 1241
verify(op === 'b00000000, "Assert 4965 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4966 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4967 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1243
#2;

verify(ir === 'b0000, "Assert 4968 : < ir !== 'b0000 >");	// Vector No: 1242
verify(op === 'b00000000, "Assert 4969 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4970 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4971 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000000100000011111100000000000000000000:1:1:0001:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000000100000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1244
#2;

verify(ir === 'b0001, "Assert 4972 : < ir !== 'b0001 >");	// Vector No: 1243
verify(op === 'b00000011, "Assert 4973 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 4974 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 4975 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000100000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000001:
//------------------------

#2;
word <= 'b0000001111110000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1245
#2;

verify(ir === 'b0000, "Assert 4976 : < ir !== 'b0000 >");	// Vector No: 1244
verify(op === 'b00000000, "Assert 4977 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4978 : < extop !== 1 >");
verify(addr === 'b00000000000000000001, "Assert 4979 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000001111110000000000000000000100000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000100000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1246
#2;

verify(ir === 'b0000, "Assert 4980 : < ir !== 'b0000 >");	// Vector No: 1245
verify(op === 'b00000000, "Assert 4981 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4982 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4983 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000100000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1247
#2;

verify(ir === 'b0011, "Assert 4984 : < ir !== 'b0011 >");	// Vector No: 1246
verify(op === 'b11110000, "Assert 4985 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 4986 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4987 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000100000000000000000000000000000000:1:1:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000100000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1248
#2;

verify(ir === 'b0001, "Assert 4988 : < ir !== 'b0001 >");	// Vector No: 1247
verify(op === 'b00000000, "Assert 4989 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4990 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 4991 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1249
#2;

verify(ir === 'b0000, "Assert 4992 : < ir !== 'b0000 >");	// Vector No: 1248
verify(op === 'b00000000, "Assert 4993 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 4994 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 4995 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1250
#2;

verify(ir === 'b0000, "Assert 4996 : < ir !== 'b0000 >");	// Vector No: 1249
verify(op === 'b00000000, "Assert 4997 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 4998 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 4999 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1251
#2;

verify(ir === 'b0000, "Assert 5000 : < ir !== 'b0000 >");	// Vector No: 1250
verify(op === 'b00000000, "Assert 5001 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5002 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5003 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000001000000011111100000000000000000000:1:1:0010:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000001000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1252
#2;

verify(ir === 'b0010, "Assert 5004 : < ir !== 'b0010 >");	// Vector No: 1251
verify(op === 'b00000011, "Assert 5005 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5006 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5007 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000001000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000010:
//------------------------

#2;
word <= 'b0000001111110000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1253
#2;

verify(ir === 'b0000, "Assert 5008 : < ir !== 'b0000 >");	// Vector No: 1252
verify(op === 'b00000000, "Assert 5009 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5010 : < extop !== 1 >");
verify(addr === 'b00000000000000000010, "Assert 5011 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000001111110000000000000000001000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000001000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1254
#2;

verify(ir === 'b0000, "Assert 5012 : < ir !== 'b0000 >");	// Vector No: 1253
verify(op === 'b00000000, "Assert 5013 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5014 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5015 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000001000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1255
#2;

verify(ir === 'b0011, "Assert 5016 : < ir !== 'b0011 >");	// Vector No: 1254
verify(op === 'b11110000, "Assert 5017 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5018 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5019 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000001000000000000000000000000000000000:1:1:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000001000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1256
#2;

verify(ir === 'b0010, "Assert 5020 : < ir !== 'b0010 >");	// Vector No: 1255
verify(op === 'b00000000, "Assert 5021 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5022 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5023 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1257
#2;

verify(ir === 'b0000, "Assert 5024 : < ir !== 'b0000 >");	// Vector No: 1256
verify(op === 'b00000000, "Assert 5025 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5026 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 5027 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1258
#2;

verify(ir === 'b0000, "Assert 5028 : < ir !== 'b0000 >");	// Vector No: 1257
verify(op === 'b00000000, "Assert 5029 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5030 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5031 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1259
#2;

verify(ir === 'b0000, "Assert 5032 : < ir !== 'b0000 >");	// Vector No: 1258
verify(op === 'b00000000, "Assert 5033 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5034 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5035 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000010000000011111100000000000000000000:1:1:0100:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000010000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1260
#2;

verify(ir === 'b0100, "Assert 5036 : < ir !== 'b0100 >");	// Vector No: 1259
verify(op === 'b00000011, "Assert 5037 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5038 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5039 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000010000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000100:
//------------------------

#2;
word <= 'b0000001111110000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1261
#2;

verify(ir === 'b0000, "Assert 5040 : < ir !== 'b0000 >");	// Vector No: 1260
verify(op === 'b00000000, "Assert 5041 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5042 : < extop !== 1 >");
verify(addr === 'b00000000000000000100, "Assert 5043 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000001111110000000000000000010000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000010000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1262
#2;

verify(ir === 'b0000, "Assert 5044 : < ir !== 'b0000 >");	// Vector No: 1261
verify(op === 'b00000000, "Assert 5045 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5046 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5047 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000010000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1263
#2;

verify(ir === 'b0011, "Assert 5048 : < ir !== 'b0011 >");	// Vector No: 1262
verify(op === 'b11110000, "Assert 5049 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5050 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5051 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000010000000000000000000000000000000000:1:1:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000010000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1264
#2;

verify(ir === 'b0100, "Assert 5052 : < ir !== 'b0100 >");	// Vector No: 1263
verify(op === 'b00000000, "Assert 5053 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5054 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5055 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1265
#2;

verify(ir === 'b0000, "Assert 5056 : < ir !== 'b0000 >");	// Vector No: 1264
verify(op === 'b00000000, "Assert 5057 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5058 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 5059 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1266
#2;

verify(ir === 'b0000, "Assert 5060 : < ir !== 'b0000 >");	// Vector No: 1265
verify(op === 'b00000000, "Assert 5061 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5062 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5063 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1267
#2;

verify(ir === 'b0000, "Assert 5064 : < ir !== 'b0000 >");	// Vector No: 1266
verify(op === 'b00000000, "Assert 5065 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5066 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5067 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000000100000000011111100000000000000000000:1:1:1000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000000100000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1268
#2;

verify(ir === 'b1000, "Assert 5068 : < ir !== 'b1000 >");	// Vector No: 1267
verify(op === 'b00000011, "Assert 5069 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5070 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5071 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000100000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000001000:
//------------------------

#2;
word <= 'b0000001111110000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1269
#2;

verify(ir === 'b0000, "Assert 5072 : < ir !== 'b0000 >");	// Vector No: 1268
verify(op === 'b00000000, "Assert 5073 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5074 : < extop !== 1 >");
verify(addr === 'b00000000000000001000, "Assert 5075 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000001111110000000000000000100000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000100000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1270
#2;

verify(ir === 'b0000, "Assert 5076 : < ir !== 'b0000 >");	// Vector No: 1269
verify(op === 'b00000000, "Assert 5077 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5078 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5079 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000100000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1271
#2;

verify(ir === 'b0011, "Assert 5080 : < ir !== 'b0011 >");	// Vector No: 1270
verify(op === 'b11110000, "Assert 5081 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5082 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5083 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000100000000000000000000000000000000000:1:1:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000100000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1272
#2;

verify(ir === 'b1000, "Assert 5084 : < ir !== 'b1000 >");	// Vector No: 1271
verify(op === 'b00000000, "Assert 5085 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5086 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5087 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1273
#2;

verify(ir === 'b0000, "Assert 5088 : < ir !== 'b0000 >");	// Vector No: 1272
verify(op === 'b00000000, "Assert 5089 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5090 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 5091 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1274
#2;

verify(ir === 'b0000, "Assert 5092 : < ir !== 'b0000 >");	// Vector No: 1273
verify(op === 'b00000000, "Assert 5093 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5094 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5095 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1275
#2;

verify(ir === 'b0000, "Assert 5096 : < ir !== 'b0000 >");	// Vector No: 1274
verify(op === 'b00000000, "Assert 5097 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5098 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 5099 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000000000000000000000000001000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000001000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1276
#2;

verify(ir === 'b0000, "Assert 5100 : < ir !== 'b0000 >");	// Vector No: 1275
verify(op === 'b00000011, "Assert 5101 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5102 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5103 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000001000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000010000:
//------------------------

#2;
word <= 'b0000001111110000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1277
#2;

verify(ir === 'b0000, "Assert 5104 : < ir !== 'b0000 >");	// Vector No: 1276
verify(op === 'b00000000, "Assert 5105 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5106 : < extop !== 1 >");
verify(addr === 'b00000000000000010000, "Assert 5107 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000001111110000000000000001000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000001000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1278
#2;

verify(ir === 'b0000, "Assert 5108 : < ir !== 'b0000 >");	// Vector No: 1277
verify(op === 'b00000000, "Assert 5109 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5110 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5111 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000001000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000001:
//------------------------

#2;
word <= 'b0000001111110000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1279
#2;

verify(ir === 'b0011, "Assert 5112 : < ir !== 'b0011 >");	// Vector No: 1278
verify(op === 'b11110000, "Assert 5113 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5114 : < extop !== 0 >");
verify(addr === 'b00000000000000000001, "Assert 5115 : < addr !== 'b00000000000000000001 >");
#2;
clk <= 0;

// 0000001111110000000000000001000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000001000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1280
#2;

verify(ir === 'b0000, "Assert 5116 : < ir !== 'b0000 >");	// Vector No: 1279
verify(op === 'b00000000, "Assert 5117 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5118 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5119 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1281
#2;

verify(ir === 'b0000, "Assert 5120 : < ir !== 'b0000 >");	// Vector No: 1280
verify(op === 'b00000000, "Assert 5121 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5122 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 5123 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1282
#2;

verify(ir === 'b0000, "Assert 5124 : < ir !== 'b0000 >");	// Vector No: 1281
verify(op === 'b00000000, "Assert 5125 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5126 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5127 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1283
#2;

verify(ir === 'b0000, "Assert 5128 : < ir !== 'b0000 >");	// Vector No: 1282
verify(op === 'b00000000, "Assert 5129 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5130 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 5131 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000000000000000000000000010000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000010000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1284
#2;

verify(ir === 'b0000, "Assert 5132 : < ir !== 'b0000 >");	// Vector No: 1283
verify(op === 'b00000011, "Assert 5133 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5134 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5135 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000010000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000100000:
//------------------------

#2;
word <= 'b0000001111110000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1285
#2;

verify(ir === 'b0000, "Assert 5136 : < ir !== 'b0000 >");	// Vector No: 1284
verify(op === 'b00000000, "Assert 5137 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5138 : < extop !== 1 >");
verify(addr === 'b00000000000000100000, "Assert 5139 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000001111110000000000000010000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000010000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1286
#2;

verify(ir === 'b0000, "Assert 5140 : < ir !== 'b0000 >");	// Vector No: 1285
verify(op === 'b00000000, "Assert 5141 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5142 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5143 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000010000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000010:
//------------------------

#2;
word <= 'b0000001111110000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1287
#2;

verify(ir === 'b0011, "Assert 5144 : < ir !== 'b0011 >");	// Vector No: 1286
verify(op === 'b11110000, "Assert 5145 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5146 : < extop !== 0 >");
verify(addr === 'b00000000000000000010, "Assert 5147 : < addr !== 'b00000000000000000010 >");
#2;
clk <= 0;

// 0000001111110000000000000010000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000010000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1288
#2;

verify(ir === 'b0000, "Assert 5148 : < ir !== 'b0000 >");	// Vector No: 1287
verify(op === 'b00000000, "Assert 5149 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5150 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5151 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1289
#2;

verify(ir === 'b0000, "Assert 5152 : < ir !== 'b0000 >");	// Vector No: 1288
verify(op === 'b00000000, "Assert 5153 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5154 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 5155 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1290
#2;

verify(ir === 'b0000, "Assert 5156 : < ir !== 'b0000 >");	// Vector No: 1289
verify(op === 'b00000000, "Assert 5157 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5158 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5159 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1291
#2;

verify(ir === 'b0000, "Assert 5160 : < ir !== 'b0000 >");	// Vector No: 1290
verify(op === 'b00000000, "Assert 5161 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5162 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 5163 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000000000000000000000000100000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000000100000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1292
#2;

verify(ir === 'b0000, "Assert 5164 : < ir !== 'b0000 >");	// Vector No: 1291
verify(op === 'b00000011, "Assert 5165 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5166 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5167 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000100000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000001000000:
//------------------------

#2;
word <= 'b0000001111110000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1293
#2;

verify(ir === 'b0000, "Assert 5168 : < ir !== 'b0000 >");	// Vector No: 1292
verify(op === 'b00000000, "Assert 5169 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5170 : < extop !== 1 >");
verify(addr === 'b00000000000001000000, "Assert 5171 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000001111110000000000000100000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000100000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1294
#2;

verify(ir === 'b0000, "Assert 5172 : < ir !== 'b0000 >");	// Vector No: 1293
verify(op === 'b00000000, "Assert 5173 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5174 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5175 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000100000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000100:
//------------------------

#2;
word <= 'b0000001111110000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1295
#2;

verify(ir === 'b0011, "Assert 5176 : < ir !== 'b0011 >");	// Vector No: 1294
verify(op === 'b11110000, "Assert 5177 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5178 : < extop !== 0 >");
verify(addr === 'b00000000000000000100, "Assert 5179 : < addr !== 'b00000000000000000100 >");
#2;
clk <= 0;

// 0000001111110000000000000100000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000100000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1296
#2;

verify(ir === 'b0000, "Assert 5180 : < ir !== 'b0000 >");	// Vector No: 1295
verify(op === 'b00000000, "Assert 5181 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5182 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5183 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1297
#2;

verify(ir === 'b0000, "Assert 5184 : < ir !== 'b0000 >");	// Vector No: 1296
verify(op === 'b00000000, "Assert 5185 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5186 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 5187 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1298
#2;

verify(ir === 'b0000, "Assert 5188 : < ir !== 'b0000 >");	// Vector No: 1297
verify(op === 'b00000000, "Assert 5189 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5190 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5191 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1299
#2;

verify(ir === 'b0000, "Assert 5192 : < ir !== 'b0000 >");	// Vector No: 1298
verify(op === 'b00000000, "Assert 5193 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5194 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 5195 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000000000000000000000001000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000001000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1300
#2;

verify(ir === 'b0000, "Assert 5196 : < ir !== 'b0000 >");	// Vector No: 1299
verify(op === 'b00000011, "Assert 5197 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5198 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5199 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000001000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000010000000:
//------------------------

#2;
word <= 'b0000001111110000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1301
#2;

verify(ir === 'b0000, "Assert 5200 : < ir !== 'b0000 >");	// Vector No: 1300
verify(op === 'b00000000, "Assert 5201 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5202 : < extop !== 1 >");
verify(addr === 'b00000000000010000000, "Assert 5203 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000001111110000000000001000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000001000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1302
#2;

verify(ir === 'b0000, "Assert 5204 : < ir !== 'b0000 >");	// Vector No: 1301
verify(op === 'b00000000, "Assert 5205 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5206 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5207 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000001000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000001000:
//------------------------

#2;
word <= 'b0000001111110000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1303
#2;

verify(ir === 'b0011, "Assert 5208 : < ir !== 'b0011 >");	// Vector No: 1302
verify(op === 'b11110000, "Assert 5209 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5210 : < extop !== 0 >");
verify(addr === 'b00000000000000001000, "Assert 5211 : < addr !== 'b00000000000000001000 >");
#2;
clk <= 0;

// 0000001111110000000000001000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000001000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1304
#2;

verify(ir === 'b0000, "Assert 5212 : < ir !== 'b0000 >");	// Vector No: 1303
verify(op === 'b00000000, "Assert 5213 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5214 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5215 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1305
#2;

verify(ir === 'b0000, "Assert 5216 : < ir !== 'b0000 >");	// Vector No: 1304
verify(op === 'b00000000, "Assert 5217 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5218 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 5219 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1306
#2;

verify(ir === 'b0000, "Assert 5220 : < ir !== 'b0000 >");	// Vector No: 1305
verify(op === 'b00000000, "Assert 5221 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5222 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5223 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1307
#2;

verify(ir === 'b0000, "Assert 5224 : < ir !== 'b0000 >");	// Vector No: 1306
verify(op === 'b00000000, "Assert 5225 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5226 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 5227 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000000000000000000000010000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000010000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1308
#2;

verify(ir === 'b0000, "Assert 5228 : < ir !== 'b0000 >");	// Vector No: 1307
verify(op === 'b00000011, "Assert 5229 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5230 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5231 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000010000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000100000000:
//------------------------

#2;
word <= 'b0000001111110000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1309
#2;

verify(ir === 'b0000, "Assert 5232 : < ir !== 'b0000 >");	// Vector No: 1308
verify(op === 'b00000000, "Assert 5233 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5234 : < extop !== 1 >");
verify(addr === 'b00000000000100000000, "Assert 5235 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000001111110000000000010000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000010000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1310
#2;

verify(ir === 'b0000, "Assert 5236 : < ir !== 'b0000 >");	// Vector No: 1309
verify(op === 'b00000000, "Assert 5237 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5238 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5239 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000010000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000010000:
//------------------------

#2;
word <= 'b0000001111110000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1311
#2;

verify(ir === 'b0011, "Assert 5240 : < ir !== 'b0011 >");	// Vector No: 1310
verify(op === 'b11110000, "Assert 5241 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5242 : < extop !== 0 >");
verify(addr === 'b00000000000000010000, "Assert 5243 : < addr !== 'b00000000000000010000 >");
#2;
clk <= 0;

// 0000001111110000000000010000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000010000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1312
#2;

verify(ir === 'b0000, "Assert 5244 : < ir !== 'b0000 >");	// Vector No: 1311
verify(op === 'b00000000, "Assert 5245 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5246 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5247 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1313
#2;

verify(ir === 'b0000, "Assert 5248 : < ir !== 'b0000 >");	// Vector No: 1312
verify(op === 'b00000000, "Assert 5249 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5250 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 5251 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1314
#2;

verify(ir === 'b0000, "Assert 5252 : < ir !== 'b0000 >");	// Vector No: 1313
verify(op === 'b00000000, "Assert 5253 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5254 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5255 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1315
#2;

verify(ir === 'b0000, "Assert 5256 : < ir !== 'b0000 >");	// Vector No: 1314
verify(op === 'b00000000, "Assert 5257 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5258 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 5259 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000000000000000000000100000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000000100000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1316
#2;

verify(ir === 'b0000, "Assert 5260 : < ir !== 'b0000 >");	// Vector No: 1315
verify(op === 'b00000011, "Assert 5261 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5262 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5263 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000100000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000001000000000:
//------------------------

#2;
word <= 'b0000001111110000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1317
#2;

verify(ir === 'b0000, "Assert 5264 : < ir !== 'b0000 >");	// Vector No: 1316
verify(op === 'b00000000, "Assert 5265 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5266 : < extop !== 1 >");
verify(addr === 'b00000000001000000000, "Assert 5267 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000001111110000000000100000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000100000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1318
#2;

verify(ir === 'b0000, "Assert 5268 : < ir !== 'b0000 >");	// Vector No: 1317
verify(op === 'b00000000, "Assert 5269 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5270 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5271 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000100000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000100000:
//------------------------

#2;
word <= 'b0000001111110000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1319
#2;

verify(ir === 'b0011, "Assert 5272 : < ir !== 'b0011 >");	// Vector No: 1318
verify(op === 'b11110000, "Assert 5273 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5274 : < extop !== 0 >");
verify(addr === 'b00000000000000100000, "Assert 5275 : < addr !== 'b00000000000000100000 >");
#2;
clk <= 0;

// 0000001111110000000000100000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000100000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1320
#2;

verify(ir === 'b0000, "Assert 5276 : < ir !== 'b0000 >");	// Vector No: 1319
verify(op === 'b00000000, "Assert 5277 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5278 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5279 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1321
#2;

verify(ir === 'b0000, "Assert 5280 : < ir !== 'b0000 >");	// Vector No: 1320
verify(op === 'b00000000, "Assert 5281 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5282 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 5283 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1322
#2;

verify(ir === 'b0000, "Assert 5284 : < ir !== 'b0000 >");	// Vector No: 1321
verify(op === 'b00000000, "Assert 5285 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5286 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5287 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1323
#2;

verify(ir === 'b0000, "Assert 5288 : < ir !== 'b0000 >");	// Vector No: 1322
verify(op === 'b00000000, "Assert 5289 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5290 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 5291 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000000000000000000001000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000001000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1324
#2;

verify(ir === 'b0000, "Assert 5292 : < ir !== 'b0000 >");	// Vector No: 1323
verify(op === 'b00000011, "Assert 5293 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5294 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5295 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000001000000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000010000000000:
//------------------------

#2;
word <= 'b0000001111110000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1325
#2;

verify(ir === 'b0000, "Assert 5296 : < ir !== 'b0000 >");	// Vector No: 1324
verify(op === 'b00000000, "Assert 5297 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5298 : < extop !== 1 >");
verify(addr === 'b00000000010000000000, "Assert 5299 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000001111110000000001000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000001000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1326
#2;

verify(ir === 'b0000, "Assert 5300 : < ir !== 'b0000 >");	// Vector No: 1325
verify(op === 'b00000000, "Assert 5301 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5302 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5303 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000001000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000001000000:
//------------------------

#2;
word <= 'b0000001111110000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1327
#2;

verify(ir === 'b0011, "Assert 5304 : < ir !== 'b0011 >");	// Vector No: 1326
verify(op === 'b11110000, "Assert 5305 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5306 : < extop !== 0 >");
verify(addr === 'b00000000000001000000, "Assert 5307 : < addr !== 'b00000000000001000000 >");
#2;
clk <= 0;

// 0000001111110000000001000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000001000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1328
#2;

verify(ir === 'b0000, "Assert 5308 : < ir !== 'b0000 >");	// Vector No: 1327
verify(op === 'b00000000, "Assert 5309 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5310 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5311 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1329
#2;

verify(ir === 'b0000, "Assert 5312 : < ir !== 'b0000 >");	// Vector No: 1328
verify(op === 'b00000000, "Assert 5313 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5314 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 5315 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1330
#2;

verify(ir === 'b0000, "Assert 5316 : < ir !== 'b0000 >");	// Vector No: 1329
verify(op === 'b00000000, "Assert 5317 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5318 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5319 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1331
#2;

verify(ir === 'b0000, "Assert 5320 : < ir !== 'b0000 >");	// Vector No: 1330
verify(op === 'b00000000, "Assert 5321 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5322 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 5323 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000000000000000000010000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000010000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1332
#2;

verify(ir === 'b0000, "Assert 5324 : < ir !== 'b0000 >");	// Vector No: 1331
verify(op === 'b00000011, "Assert 5325 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5326 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5327 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000010000000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000100000000000:
//------------------------

#2;
word <= 'b0000001111110000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1333
#2;

verify(ir === 'b0000, "Assert 5328 : < ir !== 'b0000 >");	// Vector No: 1332
verify(op === 'b00000000, "Assert 5329 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5330 : < extop !== 1 >");
verify(addr === 'b00000000100000000000, "Assert 5331 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000001111110000000010000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000010000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1334
#2;

verify(ir === 'b0000, "Assert 5332 : < ir !== 'b0000 >");	// Vector No: 1333
verify(op === 'b00000000, "Assert 5333 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5334 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5335 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000010000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000010000000:
//------------------------

#2;
word <= 'b0000001111110000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1335
#2;

verify(ir === 'b0011, "Assert 5336 : < ir !== 'b0011 >");	// Vector No: 1334
verify(op === 'b11110000, "Assert 5337 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5338 : < extop !== 0 >");
verify(addr === 'b00000000000010000000, "Assert 5339 : < addr !== 'b00000000000010000000 >");
#2;
clk <= 0;

// 0000001111110000000010000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000010000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1336
#2;

verify(ir === 'b0000, "Assert 5340 : < ir !== 'b0000 >");	// Vector No: 1335
verify(op === 'b00000000, "Assert 5341 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5342 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5343 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1337
#2;

verify(ir === 'b0000, "Assert 5344 : < ir !== 'b0000 >");	// Vector No: 1336
verify(op === 'b00000000, "Assert 5345 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5346 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 5347 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1338
#2;

verify(ir === 'b0000, "Assert 5348 : < ir !== 'b0000 >");	// Vector No: 1337
verify(op === 'b00000000, "Assert 5349 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5350 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5351 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1339
#2;

verify(ir === 'b0000, "Assert 5352 : < ir !== 'b0000 >");	// Vector No: 1338
verify(op === 'b00000000, "Assert 5353 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5354 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 5355 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000000000000000000100000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000000100000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1340
#2;

verify(ir === 'b0000, "Assert 5356 : < ir !== 'b0000 >");	// Vector No: 1339
verify(op === 'b00000011, "Assert 5357 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5358 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5359 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000100000000000000000000000000000000000000000000:0:0:0000:00000001:1:00000001000000000000:
//------------------------

#2;
word <= 'b0000001111110000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1341
#2;

verify(ir === 'b0000, "Assert 5360 : < ir !== 'b0000 >");	// Vector No: 1340
verify(op === 'b00000001, "Assert 5361 : < op !== 'b00000001 >");
verify(extop === 1, "Assert 5362 : < extop !== 1 >");
verify(addr === 'b00000001000000000000, "Assert 5363 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000001111110000000100000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000100000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1342
#2;

verify(ir === 'b0000, "Assert 5364 : < ir !== 'b0000 >");	// Vector No: 1341
verify(op === 'b00000000, "Assert 5365 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5366 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5367 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000100000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000100000000:
//------------------------

#2;
word <= 'b0000001111110000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1343
#2;

verify(ir === 'b0011, "Assert 5368 : < ir !== 'b0011 >");	// Vector No: 1342
verify(op === 'b11110000, "Assert 5369 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5370 : < extop !== 0 >");
verify(addr === 'b00000000000100000000, "Assert 5371 : < addr !== 'b00000000000100000000 >");
#2;
clk <= 0;

// 0000001111110000000100000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000100000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1344
#2;

verify(ir === 'b0000, "Assert 5372 : < ir !== 'b0000 >");	// Vector No: 1343
verify(op === 'b00000000, "Assert 5373 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5374 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5375 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1345
#2;

verify(ir === 'b0000, "Assert 5376 : < ir !== 'b0000 >");	// Vector No: 1344
verify(op === 'b00000000, "Assert 5377 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5378 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 5379 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1346
#2;

verify(ir === 'b0000, "Assert 5380 : < ir !== 'b0000 >");	// Vector No: 1345
verify(op === 'b00000000, "Assert 5381 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5382 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5383 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1347
#2;

verify(ir === 'b0000, "Assert 5384 : < ir !== 'b0000 >");	// Vector No: 1346
verify(op === 'b00000000, "Assert 5385 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5386 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 5387 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000000000000000001000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000001000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1348
#2;

verify(ir === 'b0000, "Assert 5388 : < ir !== 'b0000 >");	// Vector No: 1347
verify(op === 'b00000011, "Assert 5389 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5390 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5391 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000001000000000000000000000000000000000000000000000:0:0:0000:00000010:1:00000010000000000000:
//------------------------

#2;
word <= 'b0000001111110000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1349
#2;

verify(ir === 'b0000, "Assert 5392 : < ir !== 'b0000 >");	// Vector No: 1348
verify(op === 'b00000010, "Assert 5393 : < op !== 'b00000010 >");
verify(extop === 1, "Assert 5394 : < extop !== 1 >");
verify(addr === 'b00000010000000000000, "Assert 5395 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000001111110000001000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000001000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1350
#2;

verify(ir === 'b0000, "Assert 5396 : < ir !== 'b0000 >");	// Vector No: 1349
verify(op === 'b00000000, "Assert 5397 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5398 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5399 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000001000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000001000000000:
//------------------------

#2;
word <= 'b0000001111110000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1351
#2;

verify(ir === 'b0011, "Assert 5400 : < ir !== 'b0011 >");	// Vector No: 1350
verify(op === 'b11110000, "Assert 5401 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5402 : < extop !== 0 >");
verify(addr === 'b00000000001000000000, "Assert 5403 : < addr !== 'b00000000001000000000 >");
#2;
clk <= 0;

// 0000001111110000001000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000001000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1352
#2;

verify(ir === 'b0000, "Assert 5404 : < ir !== 'b0000 >");	// Vector No: 1351
verify(op === 'b00000000, "Assert 5405 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5406 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5407 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1353
#2;

verify(ir === 'b0000, "Assert 5408 : < ir !== 'b0000 >");	// Vector No: 1352
verify(op === 'b00000000, "Assert 5409 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5410 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 5411 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1354
#2;

verify(ir === 'b0000, "Assert 5412 : < ir !== 'b0000 >");	// Vector No: 1353
verify(op === 'b00000000, "Assert 5413 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5414 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5415 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1355
#2;

verify(ir === 'b0000, "Assert 5416 : < ir !== 'b0000 >");	// Vector No: 1354
verify(op === 'b00000000, "Assert 5417 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5418 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 5419 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000000000000000010000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000010000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1356
#2;

verify(ir === 'b0000, "Assert 5420 : < ir !== 'b0000 >");	// Vector No: 1355
verify(op === 'b00000011, "Assert 5421 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5422 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5423 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000010000000000000000000000000000000000000000000000:0:0:0000:00000100:1:00000100000000000000:
//------------------------

#2;
word <= 'b0000001111110000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1357
#2;

verify(ir === 'b0000, "Assert 5424 : < ir !== 'b0000 >");	// Vector No: 1356
verify(op === 'b00000100, "Assert 5425 : < op !== 'b00000100 >");
verify(extop === 1, "Assert 5426 : < extop !== 1 >");
verify(addr === 'b00000100000000000000, "Assert 5427 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000001111110000010000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000010000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1358
#2;

verify(ir === 'b0000, "Assert 5428 : < ir !== 'b0000 >");	// Vector No: 1357
verify(op === 'b00000000, "Assert 5429 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5430 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5431 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000010000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000010000000000:
//------------------------

#2;
word <= 'b0000001111110000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1359
#2;

verify(ir === 'b0011, "Assert 5432 : < ir !== 'b0011 >");	// Vector No: 1358
verify(op === 'b11110000, "Assert 5433 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5434 : < extop !== 0 >");
verify(addr === 'b00000000010000000000, "Assert 5435 : < addr !== 'b00000000010000000000 >");
#2;
clk <= 0;

// 0000001111110000010000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000010000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1360
#2;

verify(ir === 'b0000, "Assert 5436 : < ir !== 'b0000 >");	// Vector No: 1359
verify(op === 'b00000000, "Assert 5437 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5438 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5439 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00001000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1361
#2;

verify(ir === 'b0000, "Assert 5440 : < ir !== 'b0000 >");	// Vector No: 1360
verify(op === 'b00000000, "Assert 5441 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5442 : < extop !== 0 >");
verify(addr === 'b00001000000000000000, "Assert 5443 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1362
#2;

verify(ir === 'b0000, "Assert 5444 : < ir !== 'b0000 >");	// Vector No: 1361
verify(op === 'b00000000, "Assert 5445 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5446 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5447 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1363
#2;

verify(ir === 'b0000, "Assert 5448 : < ir !== 'b0000 >");	// Vector No: 1362
verify(op === 'b00000000, "Assert 5449 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5450 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 5451 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000000000000000100000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000000100000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1364
#2;

verify(ir === 'b0000, "Assert 5452 : < ir !== 'b0000 >");	// Vector No: 1363
verify(op === 'b00000011, "Assert 5453 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5454 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5455 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000100000000000000000000000000000000000000000000000:0:0:0000:00001000:1:00001000000000000000:
//------------------------

#2;
word <= 'b0000001111110000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1365
#2;

verify(ir === 'b0000, "Assert 5456 : < ir !== 'b0000 >");	// Vector No: 1364
verify(op === 'b00001000, "Assert 5457 : < op !== 'b00001000 >");
verify(extop === 1, "Assert 5458 : < extop !== 1 >");
verify(addr === 'b00001000000000000000, "Assert 5459 : < addr !== 'b00001000000000000000 >");
#2;
clk <= 0;

// 0000001111110000100000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000100000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1366
#2;

verify(ir === 'b0000, "Assert 5460 : < ir !== 'b0000 >");	// Vector No: 1365
verify(op === 'b00000000, "Assert 5461 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5462 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5463 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000100000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000100000000000:
//------------------------

#2;
word <= 'b0000001111110000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1367
#2;

verify(ir === 'b0011, "Assert 5464 : < ir !== 'b0011 >");	// Vector No: 1366
verify(op === 'b11110000, "Assert 5465 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5466 : < extop !== 0 >");
verify(addr === 'b00000000100000000000, "Assert 5467 : < addr !== 'b00000000100000000000 >");
#2;
clk <= 0;

// 0000001111110000100000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000100000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1368
#2;

verify(ir === 'b0000, "Assert 5468 : < ir !== 'b0000 >");	// Vector No: 1367
verify(op === 'b00000000, "Assert 5469 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5470 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5471 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00010000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1369
#2;

verify(ir === 'b0000, "Assert 5472 : < ir !== 'b0000 >");	// Vector No: 1368
verify(op === 'b00000000, "Assert 5473 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5474 : < extop !== 0 >");
verify(addr === 'b00010000000000000000, "Assert 5475 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1370
#2;

verify(ir === 'b0000, "Assert 5476 : < ir !== 'b0000 >");	// Vector No: 1369
verify(op === 'b00000000, "Assert 5477 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5478 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5479 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000011111100000000000000000000:1:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1371
#2;

verify(ir === 'b0000, "Assert 5480 : < ir !== 'b0000 >");	// Vector No: 1370
verify(op === 'b00000001, "Assert 5481 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 5482 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5483 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000001000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000001000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1372
#2;

verify(ir === 'b0000, "Assert 5484 : < ir !== 'b0000 >");	// Vector No: 1371
verify(op === 'b00000011, "Assert 5485 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5486 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5487 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110001000000000000000000000000000000000000000000000000:0:0:0000:00010000:1:00010000000000000000:
//------------------------

#2;
word <= 'b0000001111110001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1373
#2;

verify(ir === 'b0000, "Assert 5488 : < ir !== 'b0000 >");	// Vector No: 1372
verify(op === 'b00010000, "Assert 5489 : < op !== 'b00010000 >");
verify(extop === 1, "Assert 5490 : < extop !== 1 >");
verify(addr === 'b00010000000000000000, "Assert 5491 : < addr !== 'b00010000000000000000 >");
#2;
clk <= 0;

// 0000001111110001000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110001000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1374
#2;

verify(ir === 'b0000, "Assert 5492 : < ir !== 'b0000 >");	// Vector No: 1373
verify(op === 'b00000000, "Assert 5493 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5494 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5495 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110001000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000001000000000000:
//------------------------

#2;
word <= 'b0000001111110001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1375
#2;

verify(ir === 'b0011, "Assert 5496 : < ir !== 'b0011 >");	// Vector No: 1374
verify(op === 'b11110000, "Assert 5497 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5498 : < extop !== 0 >");
verify(addr === 'b00000001000000000000, "Assert 5499 : < addr !== 'b00000001000000000000 >");
#2;
clk <= 0;

// 0000001111110001000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110001000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1376
#2;

verify(ir === 'b0000, "Assert 5500 : < ir !== 'b0000 >");	// Vector No: 1375
verify(op === 'b00000000, "Assert 5501 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5502 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5503 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000011111100000000000000000000:0:0:0000:00000000:0:00100000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1377
#2;

verify(ir === 'b0000, "Assert 5504 : < ir !== 'b0000 >");	// Vector No: 1376
verify(op === 'b00000000, "Assert 5505 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5506 : < extop !== 0 >");
verify(addr === 'b00100000000000000000, "Assert 5507 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1378
#2;

verify(ir === 'b0000, "Assert 5508 : < ir !== 'b0000 >");	// Vector No: 1377
verify(op === 'b00000000, "Assert 5509 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5510 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5511 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000011111100000000000000000000:1:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1379
#2;

verify(ir === 'b0000, "Assert 5512 : < ir !== 'b0000 >");	// Vector No: 1378
verify(op === 'b00000010, "Assert 5513 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 5514 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5515 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000010000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000010000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1380
#2;

verify(ir === 'b0000, "Assert 5516 : < ir !== 'b0000 >");	// Vector No: 1379
verify(op === 'b00000011, "Assert 5517 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5518 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5519 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110010000000000000000000000000000000000000000000000000:0:0:0000:00100000:1:00100000000000000000:
//------------------------

#2;
word <= 'b0000001111110010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1381
#2;

verify(ir === 'b0000, "Assert 5520 : < ir !== 'b0000 >");	// Vector No: 1380
verify(op === 'b00100000, "Assert 5521 : < op !== 'b00100000 >");
verify(extop === 1, "Assert 5522 : < extop !== 1 >");
verify(addr === 'b00100000000000000000, "Assert 5523 : < addr !== 'b00100000000000000000 >");
#2;
clk <= 0;

// 0000001111110010000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110010000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1382
#2;

verify(ir === 'b0000, "Assert 5524 : < ir !== 'b0000 >");	// Vector No: 1381
verify(op === 'b00000000, "Assert 5525 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5526 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5527 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110010000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000010000000000000:
//------------------------

#2;
word <= 'b0000001111110010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1383
#2;

verify(ir === 'b0011, "Assert 5528 : < ir !== 'b0011 >");	// Vector No: 1382
verify(op === 'b11110000, "Assert 5529 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5530 : < extop !== 0 >");
verify(addr === 'b00000010000000000000, "Assert 5531 : < addr !== 'b00000010000000000000 >");
#2;
clk <= 0;

// 0000001111110010000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110010000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1384
#2;

verify(ir === 'b0000, "Assert 5532 : < ir !== 'b0000 >");	// Vector No: 1383
verify(op === 'b00000000, "Assert 5533 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5534 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5535 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000011111100000000000000000000:0:0:0000:00000000:0:01000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1385
#2;

verify(ir === 'b0000, "Assert 5536 : < ir !== 'b0000 >");	// Vector No: 1384
verify(op === 'b00000000, "Assert 5537 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5538 : < extop !== 0 >");
verify(addr === 'b01000000000000000000, "Assert 5539 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1386
#2;

verify(ir === 'b0000, "Assert 5540 : < ir !== 'b0000 >");	// Vector No: 1385
verify(op === 'b00000000, "Assert 5541 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5542 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5543 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000011111100000000000000000000:1:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1387
#2;

verify(ir === 'b0000, "Assert 5544 : < ir !== 'b0000 >");	// Vector No: 1386
verify(op === 'b00000100, "Assert 5545 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 5546 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5547 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000000100000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000000100000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1388
#2;

verify(ir === 'b0000, "Assert 5548 : < ir !== 'b0000 >");	// Vector No: 1387
verify(op === 'b00000011, "Assert 5549 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5550 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5551 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110100000000000000000000000000000000000000000000000000:0:0:0000:01000000:1:01000000000000000000:
//------------------------

#2;
word <= 'b0000001111110100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1389
#2;

verify(ir === 'b0000, "Assert 5552 : < ir !== 'b0000 >");	// Vector No: 1388
verify(op === 'b01000000, "Assert 5553 : < op !== 'b01000000 >");
verify(extop === 1, "Assert 5554 : < extop !== 1 >");
verify(addr === 'b01000000000000000000, "Assert 5555 : < addr !== 'b01000000000000000000 >");
#2;
clk <= 0;

// 0000001111110100000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110100000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1390
#2;

verify(ir === 'b0000, "Assert 5556 : < ir !== 'b0000 >");	// Vector No: 1389
verify(op === 'b00000000, "Assert 5557 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5558 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5559 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110100000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000100000000000000:
//------------------------

#2;
word <= 'b0000001111110100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1391
#2;

verify(ir === 'b0011, "Assert 5560 : < ir !== 'b0011 >");	// Vector No: 1390
verify(op === 'b11110000, "Assert 5561 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5562 : < extop !== 0 >");
verify(addr === 'b00000100000000000000, "Assert 5563 : < addr !== 'b00000100000000000000 >");
#2;
clk <= 0;

// 0000001111110100000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110100000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1392
#2;

verify(ir === 'b0000, "Assert 5564 : < ir !== 'b0000 >");	// Vector No: 1391
verify(op === 'b00000000, "Assert 5565 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5566 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5567 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000011111100000000000000000000:0:0:0000:00000000:0:10000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1393
#2;

verify(ir === 'b0000, "Assert 5568 : < ir !== 'b0000 >");	// Vector No: 1392
verify(op === 'b00000000, "Assert 5569 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5570 : < extop !== 0 >");
verify(addr === 'b10000000000000000000, "Assert 5571 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1394
#2;

verify(ir === 'b0000, "Assert 5572 : < ir !== 'b0000 >");	// Vector No: 1393
verify(op === 'b00000000, "Assert 5573 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5574 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5575 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000011111100000000000000000000:1:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1395
#2;

verify(ir === 'b0000, "Assert 5576 : < ir !== 'b0000 >");	// Vector No: 1394
verify(op === 'b00001000, "Assert 5577 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 5578 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5579 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000001000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000001000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1396
#2;

verify(ir === 'b0000, "Assert 5580 : < ir !== 'b0000 >");	// Vector No: 1395
verify(op === 'b00000011, "Assert 5581 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5582 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5583 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111111000000000000000000000000000000000000000000000000000:0:0:0000:10000000:1:10000000000000000000:
//------------------------

#2;
word <= 'b0000001111111000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1397
#2;

verify(ir === 'b0000, "Assert 5584 : < ir !== 'b0000 >");	// Vector No: 1396
verify(op === 'b10000000, "Assert 5585 : < op !== 'b10000000 >");
verify(extop === 1, "Assert 5586 : < extop !== 1 >");
verify(addr === 'b10000000000000000000, "Assert 5587 : < addr !== 'b10000000000000000000 >");
#2;
clk <= 0;

// 0000001111111000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111111000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1398
#2;

verify(ir === 'b0000, "Assert 5588 : < ir !== 'b0000 >");	// Vector No: 1397
verify(op === 'b00000000, "Assert 5589 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5590 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5591 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111111000000000000000000000000000000000000000000000000000:1:0:0011:11111000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111111000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1399
#2;

verify(ir === 'b0011, "Assert 5592 : < ir !== 'b0011 >");	// Vector No: 1398
verify(op === 'b11111000, "Assert 5593 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5594 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5595 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111111000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111111000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1400
#2;

verify(ir === 'b0000, "Assert 5596 : < ir !== 'b0000 >");	// Vector No: 1399
verify(op === 'b00000000, "Assert 5597 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5598 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5599 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000011111100000000000000000000:0:0:0000:00000001:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1401
#2;

verify(ir === 'b0000, "Assert 5600 : < ir !== 'b0000 >");	// Vector No: 1400
verify(op === 'b00000001, "Assert 5601 : < op !== 'b00000001 >");
verify(extop === 0, "Assert 5602 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5603 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1402
#2;

verify(ir === 'b0000, "Assert 5604 : < ir !== 'b0000 >");	// Vector No: 1401
verify(op === 'b00000000, "Assert 5605 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5606 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5607 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000011111100000000000000000000:1:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1403
#2;

verify(ir === 'b0000, "Assert 5608 : < ir !== 'b0000 >");	// Vector No: 1402
verify(op === 'b00010000, "Assert 5609 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 5610 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5611 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000010000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000010000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1404
#2;

verify(ir === 'b0000, "Assert 5612 : < ir !== 'b0000 >");	// Vector No: 1403
verify(op === 'b00000011, "Assert 5613 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5614 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5615 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000000:0:0:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1405
#2;

verify(ir === 'b0000, "Assert 5616 : < ir !== 'b0000 >");	// Vector No: 1404
verify(op === 'b00000000, "Assert 5617 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5618 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5619 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1406
#2;

verify(ir === 'b0000, "Assert 5620 : < ir !== 'b0000 >");	// Vector No: 1405
verify(op === 'b00000000, "Assert 5621 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5622 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5623 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1407
#2;

verify(ir === 'b0011, "Assert 5624 : < ir !== 'b0011 >");	// Vector No: 1406
verify(op === 'b11110000, "Assert 5625 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5626 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5627 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001111110000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1408
#2;

verify(ir === 'b0000, "Assert 5628 : < ir !== 'b0000 >");	// Vector No: 1407
verify(op === 'b00000000, "Assert 5629 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5630 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5631 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000011111100000000000000000000:0:0:0000:00000010:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1409
#2;

verify(ir === 'b0000, "Assert 5632 : < ir !== 'b0000 >");	// Vector No: 1408
verify(op === 'b00000010, "Assert 5633 : < op !== 'b00000010 >");
verify(extop === 0, "Assert 5634 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5635 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1410
#2;

verify(ir === 'b0000, "Assert 5636 : < ir !== 'b0000 >");	// Vector No: 1409
verify(op === 'b00000000, "Assert 5637 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5638 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5639 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000011111100000000000000000000:1:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1411
#2;

verify(ir === 'b0000, "Assert 5640 : < ir !== 'b0000 >");	// Vector No: 1410
verify(op === 'b00100000, "Assert 5641 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 5642 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5643 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000000100000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000000100000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1412
#2;

verify(ir === 'b0000, "Assert 5644 : < ir !== 'b0000 >");	// Vector No: 1411
verify(op === 'b00000011, "Assert 5645 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5646 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5647 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000011111100000000000000000000:0:0:0000:00000100:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1413
#2;

verify(ir === 'b0000, "Assert 5648 : < ir !== 'b0000 >");	// Vector No: 1412
verify(op === 'b00000100, "Assert 5649 : < op !== 'b00000100 >");
verify(extop === 0, "Assert 5650 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5651 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1414
#2;

verify(ir === 'b0000, "Assert 5652 : < ir !== 'b0000 >");	// Vector No: 1413
verify(op === 'b00000000, "Assert 5653 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5654 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5655 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000011111100000000000000000000:1:0:0000:01000000:0:00000111000000000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1415
#2;

verify(ir === 'b0000, "Assert 5656 : < ir !== 'b0000 >");	// Vector No: 1414
verify(op === 'b01000000, "Assert 5657 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 5658 : < extop !== 0 >");
verify(addr === 'b00000111000000000000, "Assert 5659 : < addr !== 'b00000111000000000000 >");
#2;
clk <= 0;

// 0000000001000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000001000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1416
#2;

verify(ir === 'b0000, "Assert 5660 : < ir !== 'b0000 >");	// Vector No: 1415
verify(op === 'b00000011, "Assert 5661 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5662 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5663 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000011111100000000000000000000:0:0:0000:00001000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1417
#2;

verify(ir === 'b0000, "Assert 5664 : < ir !== 'b0000 >");	// Vector No: 1416
verify(op === 'b00001000, "Assert 5665 : < op !== 'b00001000 >");
verify(extop === 0, "Assert 5666 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5667 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1418
#2;

verify(ir === 'b0000, "Assert 5668 : < ir !== 'b0000 >");	// Vector No: 1417
verify(op === 'b00000000, "Assert 5669 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5670 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5671 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000011111100000000000000000000:1:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1419
#2;

verify(ir === 'b0000, "Assert 5672 : < ir !== 'b0000 >");	// Vector No: 1418
verify(op === 'b10000000, "Assert 5673 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 5674 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5675 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000010000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000010000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1420
#2;

verify(ir === 'b0000, "Assert 5676 : < ir !== 'b0000 >");	// Vector No: 1419
verify(op === 'b00000011, "Assert 5677 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5678 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5679 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000011111100000000000000000000:0:0:0000:00010000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1421
#2;

verify(ir === 'b0000, "Assert 5680 : < ir !== 'b0000 >");	// Vector No: 1420
verify(op === 'b00010000, "Assert 5681 : < op !== 'b00010000 >");
verify(extop === 0, "Assert 5682 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5683 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1422
#2;

verify(ir === 'b0000, "Assert 5684 : < ir !== 'b0000 >");	// Vector No: 1421
verify(op === 'b00000000, "Assert 5685 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5686 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5687 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000011111100000000000000000000:1:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1423
#2;

verify(ir === 'b0001, "Assert 5688 : < ir !== 'b0001 >");	// Vector No: 1422
verify(op === 'b00000000, "Assert 5689 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5690 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5691 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000000100000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000000100000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1424
#2;

verify(ir === 'b0000, "Assert 5692 : < ir !== 'b0000 >");	// Vector No: 1423
verify(op === 'b00000011, "Assert 5693 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5694 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5695 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000011111100000000000000000000:0:0:0000:00100000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1425
#2;

verify(ir === 'b0000, "Assert 5696 : < ir !== 'b0000 >");	// Vector No: 1424
verify(op === 'b00100000, "Assert 5697 : < op !== 'b00100000 >");
verify(extop === 0, "Assert 5698 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5699 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1426
#2;

verify(ir === 'b0000, "Assert 5700 : < ir !== 'b0000 >");	// Vector No: 1425
verify(op === 'b00000000, "Assert 5701 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5702 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5703 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000011111100000000000000000000:1:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1427
#2;

verify(ir === 'b0010, "Assert 5704 : < ir !== 'b0010 >");	// Vector No: 1426
verify(op === 'b00000000, "Assert 5705 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5706 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5707 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000001000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000001000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1428
#2;

verify(ir === 'b0000, "Assert 5708 : < ir !== 'b0000 >");	// Vector No: 1427
verify(op === 'b00000011, "Assert 5709 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5710 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5711 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000011111100000000000000000000:0:0:0000:01000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1429
#2;

verify(ir === 'b0000, "Assert 5712 : < ir !== 'b0000 >");	// Vector No: 1428
verify(op === 'b01000000, "Assert 5713 : < op !== 'b01000000 >");
verify(extop === 0, "Assert 5714 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5715 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1430
#2;

verify(ir === 'b0000, "Assert 5716 : < ir !== 'b0000 >");	// Vector No: 1429
verify(op === 'b00000000, "Assert 5717 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5718 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5719 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000011111100000000000000000000:1:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1431
#2;

verify(ir === 'b0100, "Assert 5720 : < ir !== 'b0100 >");	// Vector No: 1430
verify(op === 'b00000000, "Assert 5721 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5722 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5723 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000010000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000010000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1432
#2;

verify(ir === 'b0000, "Assert 5724 : < ir !== 'b0000 >");	// Vector No: 1431
verify(op === 'b00000011, "Assert 5725 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5726 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5727 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000011111100000000000000000000:0:0:0000:10000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1433
#2;

verify(ir === 'b0000, "Assert 5728 : < ir !== 'b0000 >");	// Vector No: 1432
verify(op === 'b10000000, "Assert 5729 : < op !== 'b10000000 >");
verify(extop === 0, "Assert 5730 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5731 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1434
#2;

verify(ir === 'b0000, "Assert 5732 : < ir !== 'b0000 >");	// Vector No: 1433
verify(op === 'b00000000, "Assert 5733 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5734 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5735 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1435
#2;

verify(ir === 'b0000, "Assert 5736 : < ir !== 'b0000 >");	// Vector No: 1434
verify(op === 'b00000000, "Assert 5737 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5738 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5739 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0000100000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0000100000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1436
#2;

verify(ir === 'b0000, "Assert 5740 : < ir !== 'b0000 >");	// Vector No: 1435
verify(op === 'b00000011, "Assert 5741 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5742 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5743 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000011111100000000000000000000:0:0:0001:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1437
#2;

verify(ir === 'b0001, "Assert 5744 : < ir !== 'b0001 >");	// Vector No: 1436
verify(op === 'b00000000, "Assert 5745 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5746 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5747 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1438
#2;

verify(ir === 'b0000, "Assert 5748 : < ir !== 'b0000 >");	// Vector No: 1437
verify(op === 'b00000000, "Assert 5749 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5750 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5751 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1439
#2;

verify(ir === 'b0000, "Assert 5752 : < ir !== 'b0000 >");	// Vector No: 1438
verify(op === 'b00000000, "Assert 5753 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5754 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5755 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001000000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0001000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1440
#2;

verify(ir === 'b0000, "Assert 5756 : < ir !== 'b0000 >");	// Vector No: 1439
verify(op === 'b00000011, "Assert 5757 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5758 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5759 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0001001111110000000000000000000000000000000000000000000000000000:0:0:0001:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0001001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1441
#2;

verify(ir === 'b0001, "Assert 5760 : < ir !== 'b0001 >");	// Vector No: 1440
verify(op === 'b00000000, "Assert 5761 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5762 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5763 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001001111110000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1442
#2;

verify(ir === 'b0000, "Assert 5764 : < ir !== 'b0000 >");	// Vector No: 1441
verify(op === 'b00000000, "Assert 5765 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5766 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5767 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001001111110000000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1443
#2;

verify(ir === 'b0011, "Assert 5768 : < ir !== 'b0011 >");	// Vector No: 1442
verify(op === 'b11110000, "Assert 5769 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5770 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5771 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0001001111110000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0001001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1444
#2;

verify(ir === 'b0000, "Assert 5772 : < ir !== 'b0000 >");	// Vector No: 1443
verify(op === 'b00000000, "Assert 5773 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5774 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5775 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000011111100000000000000000000:0:0:0010:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1445
#2;

verify(ir === 'b0010, "Assert 5776 : < ir !== 'b0010 >");	// Vector No: 1444
verify(op === 'b00000000, "Assert 5777 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5778 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5779 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1446
#2;

verify(ir === 'b0000, "Assert 5780 : < ir !== 'b0000 >");	// Vector No: 1445
verify(op === 'b00000000, "Assert 5781 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5782 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5783 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1447
#2;

verify(ir === 'b0000, "Assert 5784 : < ir !== 'b0000 >");	// Vector No: 1446
verify(op === 'b00000000, "Assert 5785 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5786 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5787 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010000000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0010000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1448
#2;

verify(ir === 'b0000, "Assert 5788 : < ir !== 'b0000 >");	// Vector No: 1447
verify(op === 'b00000011, "Assert 5789 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5790 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5791 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0010001111110000000000000000000000000000000000000000000000000000:0:0:0010:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0010001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1449
#2;

verify(ir === 'b0010, "Assert 5792 : < ir !== 'b0010 >");	// Vector No: 1448
verify(op === 'b00000000, "Assert 5793 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5794 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5795 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010001111110000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1450
#2;

verify(ir === 'b0000, "Assert 5796 : < ir !== 'b0000 >");	// Vector No: 1449
verify(op === 'b00000000, "Assert 5797 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5798 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5799 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010001111110000000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1451
#2;

verify(ir === 'b0011, "Assert 5800 : < ir !== 'b0011 >");	// Vector No: 1450
verify(op === 'b11110000, "Assert 5801 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5802 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5803 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0010001111110000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0010001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1452
#2;

verify(ir === 'b0000, "Assert 5804 : < ir !== 'b0000 >");	// Vector No: 1451
verify(op === 'b00000000, "Assert 5805 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5806 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5807 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000011111100000000000000000000:0:0:0100:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1453
#2;

verify(ir === 'b0100, "Assert 5808 : < ir !== 'b0100 >");	// Vector No: 1452
verify(op === 'b00000000, "Assert 5809 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5810 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5811 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1454
#2;

verify(ir === 'b0000, "Assert 5812 : < ir !== 'b0000 >");	// Vector No: 1453
verify(op === 'b00000000, "Assert 5813 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5814 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5815 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000011111100000000000000000000:1:0:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1455
#2;

verify(ir === 'b0000, "Assert 5816 : < ir !== 'b0000 >");	// Vector No: 1454
verify(op === 'b00000000, "Assert 5817 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5818 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5819 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100000000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b0100000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1456
#2;

verify(ir === 'b0000, "Assert 5820 : < ir !== 'b0000 >");	// Vector No: 1455
verify(op === 'b00000011, "Assert 5821 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5822 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5823 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 0100001111110000000000000000000000000000000000000000000000000000:0:0:0100:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b0100001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1457
#2;

verify(ir === 'b0100, "Assert 5824 : < ir !== 'b0100 >");	// Vector No: 1456
verify(op === 'b00000000, "Assert 5825 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5826 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5827 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100001111110000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1458
#2;

verify(ir === 'b0000, "Assert 5828 : < ir !== 'b0000 >");	// Vector No: 1457
verify(op === 'b00000000, "Assert 5829 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5830 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5831 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100001111110000000000000000000000000000000000000000000000000000:1:0:0011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1459
#2;

verify(ir === 'b0011, "Assert 5832 : < ir !== 'b0011 >");	// Vector No: 1458
verify(op === 'b11110000, "Assert 5833 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5834 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5835 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 0100001111110000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b0100001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1460
#2;

verify(ir === 'b0000, "Assert 5836 : < ir !== 'b0000 >");	// Vector No: 1459
verify(op === 'b00000000, "Assert 5837 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5838 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5839 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000011111100000000000000000000:0:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1461
#2;

verify(ir === 'b1000, "Assert 5840 : < ir !== 'b1000 >");	// Vector No: 1460
verify(op === 'b00000000, "Assert 5841 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5842 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5843 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000011111100000000000000000000:0:1:0000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000011111100000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1462
#2;

verify(ir === 'b0000, "Assert 5844 : < ir !== 'b0000 >");	// Vector No: 1461
verify(op === 'b00000000, "Assert 5845 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5846 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5847 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000011111100000000000000000000:1:0:1000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1463
#2;

verify(ir === 'b1000, "Assert 5848 : < ir !== 'b1000 >");	// Vector No: 1462
verify(op === 'b00000000, "Assert 5849 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5850 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5851 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000000000000000000000000000000000000011111100000000000000000000:1:1:0000:00000011:0:00000000111100000000:
//------------------------

#2;
word <= 'b1000000000000000000000000000000000000011111100000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1464
#2;

verify(ir === 'b0000, "Assert 5852 : < ir !== 'b0000 >");	// Vector No: 1463
verify(op === 'b00000011, "Assert 5853 : < op !== 'b00000011 >");
verify(extop === 0, "Assert 5854 : < extop !== 0 >");
verify(addr === 'b00000000111100000000, "Assert 5855 : < addr !== 'b00000000111100000000 >");
#2;
clk <= 0;

// 1000001111110000000000000000000000000000000000000000000000000000:0:0:1000:00000000:1:00000000000000000000:
//------------------------

#2;
word <= 'b1000001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1465
#2;

verify(ir === 'b1000, "Assert 5856 : < ir !== 'b1000 >");	// Vector No: 1464
verify(op === 'b00000000, "Assert 5857 : < op !== 'b00000000 >");
verify(extop === 1, "Assert 5858 : < extop !== 1 >");
verify(addr === 'b00000000000000000000, "Assert 5859 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000001111110000000000000000000000000000000000000000000000000000:0:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000001111110000000000000000000000000000000000000000000000000000;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1466
#2;

verify(ir === 'b0000, "Assert 5860 : < ir !== 'b0000 >");	// Vector No: 1465
verify(op === 'b00000000, "Assert 5861 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5862 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5863 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000001111110000000000000000000000000000000000000000000000000000:1:0:1011:11110000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1467
#2;

verify(ir === 'b1011, "Assert 5864 : < ir !== 'b1011 >");	// Vector No: 1466
verify(op === 'b11110000, "Assert 5865 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 5866 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5867 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1000001111110000000000000000000000000000000000000000000000000000:1:1:0000:00000000:0:00000000000000000000:
//------------------------

#2;
word <= 'b1000001111110000000000000000000000000000000000000000000000000000;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1468
#2;

verify(ir === 'b0000, "Assert 5868 : < ir !== 'b0000 >");	// Vector No: 1467
verify(op === 'b00000000, "Assert 5869 : < op !== 'b00000000 >");
verify(extop === 0, "Assert 5870 : < extop !== 0 >");
verify(addr === 'b00000000000000000000, "Assert 5871 : < addr !== 'b00000000000000000000 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111110:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111110;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1469
#2;

verify(ir === 'b1111, "Assert 5872 : < ir !== 'b1111 >");	// Vector No: 1468
verify(op === 'b11111111, "Assert 5873 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5874 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 5875 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111110:0:1:1111:11111111:1:11111111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111110;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1470
#2;

verify(ir === 'b1111, "Assert 5876 : < ir !== 'b1111 >");	// Vector No: 1469
verify(op === 'b11111111, "Assert 5877 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5878 : < extop !== 1 >");
verify(addr === 'b11111111111111111110, "Assert 5879 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111110:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111110;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1471
#2;

verify(ir === 'b1111, "Assert 5880 : < ir !== 'b1111 >");	// Vector No: 1470
verify(op === 'b11111000, "Assert 5881 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5882 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5883 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111110:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111110;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1472
#2;

verify(ir === 'b1111, "Assert 5884 : < ir !== 'b1111 >");	// Vector No: 1471
verify(op === 'b11100000, "Assert 5885 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 5886 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 5887 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111110:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111110;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1473
#2;

verify(ir === 'b1111, "Assert 5888 : < ir !== 'b1111 >");	// Vector No: 1472
verify(op === 'b11111111, "Assert 5889 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5890 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 5891 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111110:0:1:1111:11111111:0:11111111111111111110:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111110;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1474
#2;

verify(ir === 'b1111, "Assert 5892 : < ir !== 'b1111 >");	// Vector No: 1473
verify(op === 'b11111111, "Assert 5893 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5894 : < extop !== 0 >");
verify(addr === 'b11111111111111111110, "Assert 5895 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111110:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111110;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1475
#2;

verify(ir === 'b1011, "Assert 5896 : < ir !== 'b1011 >");	// Vector No: 1474
verify(op === 'b11111000, "Assert 5897 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5898 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5899 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111110:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111110;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1476
#2;

verify(ir === 'b1111, "Assert 5900 : < ir !== 'b1111 >");	// Vector No: 1475
verify(op === 'b11111000, "Assert 5901 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5902 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5903 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111101:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111101;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1477
#2;

verify(ir === 'b1111, "Assert 5904 : < ir !== 'b1111 >");	// Vector No: 1476
verify(op === 'b11111111, "Assert 5905 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5906 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 5907 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111101:0:1:1111:11111111:1:11111111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111101;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1478
#2;

verify(ir === 'b1111, "Assert 5908 : < ir !== 'b1111 >");	// Vector No: 1477
verify(op === 'b11111111, "Assert 5909 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5910 : < extop !== 1 >");
verify(addr === 'b11111111111111111101, "Assert 5911 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111101:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111101;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1479
#2;

verify(ir === 'b1111, "Assert 5912 : < ir !== 'b1111 >");	// Vector No: 1478
verify(op === 'b11111000, "Assert 5913 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5914 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5915 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111101:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111101;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1480
#2;

verify(ir === 'b1111, "Assert 5916 : < ir !== 'b1111 >");	// Vector No: 1479
verify(op === 'b11100000, "Assert 5917 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 5918 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 5919 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111101:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111101;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1481
#2;

verify(ir === 'b1111, "Assert 5920 : < ir !== 'b1111 >");	// Vector No: 1480
verify(op === 'b11111111, "Assert 5921 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5922 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 5923 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111101:0:1:1111:11111111:0:11111111111111111101:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111101;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1482
#2;

verify(ir === 'b1111, "Assert 5924 : < ir !== 'b1111 >");	// Vector No: 1481
verify(op === 'b11111111, "Assert 5925 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5926 : < extop !== 0 >");
verify(addr === 'b11111111111111111101, "Assert 5927 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111101:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111101;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1483
#2;

verify(ir === 'b1011, "Assert 5928 : < ir !== 'b1011 >");	// Vector No: 1482
verify(op === 'b11111000, "Assert 5929 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5930 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5931 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111101:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111101;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1484
#2;

verify(ir === 'b1111, "Assert 5932 : < ir !== 'b1111 >");	// Vector No: 1483
verify(op === 'b11111000, "Assert 5933 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5934 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5935 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111011:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111011;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1485
#2;

verify(ir === 'b1111, "Assert 5936 : < ir !== 'b1111 >");	// Vector No: 1484
verify(op === 'b11111111, "Assert 5937 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5938 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 5939 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111011:0:1:1111:11111111:1:11111111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111011;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1486
#2;

verify(ir === 'b1111, "Assert 5940 : < ir !== 'b1111 >");	// Vector No: 1485
verify(op === 'b11111111, "Assert 5941 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5942 : < extop !== 1 >");
verify(addr === 'b11111111111111111011, "Assert 5943 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111011:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111011;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1487
#2;

verify(ir === 'b1111, "Assert 5944 : < ir !== 'b1111 >");	// Vector No: 1486
verify(op === 'b11111000, "Assert 5945 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5946 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5947 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111011:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111011;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1488
#2;

verify(ir === 'b1111, "Assert 5948 : < ir !== 'b1111 >");	// Vector No: 1487
verify(op === 'b11100000, "Assert 5949 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 5950 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 5951 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111011:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111011;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1489
#2;

verify(ir === 'b1111, "Assert 5952 : < ir !== 'b1111 >");	// Vector No: 1488
verify(op === 'b11111111, "Assert 5953 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5954 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 5955 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111011:0:1:1111:11111111:0:11111111111111111011:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111011;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1490
#2;

verify(ir === 'b1111, "Assert 5956 : < ir !== 'b1111 >");	// Vector No: 1489
verify(op === 'b11111111, "Assert 5957 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5958 : < extop !== 0 >");
verify(addr === 'b11111111111111111011, "Assert 5959 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111011:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111011;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1491
#2;

verify(ir === 'b1011, "Assert 5960 : < ir !== 'b1011 >");	// Vector No: 1490
verify(op === 'b11111000, "Assert 5961 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5962 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5963 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111011:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111011;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1492
#2;

verify(ir === 'b1111, "Assert 5964 : < ir !== 'b1111 >");	// Vector No: 1491
verify(op === 'b11111000, "Assert 5965 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5966 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5967 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111110111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111110111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1493
#2;

verify(ir === 'b1111, "Assert 5968 : < ir !== 'b1111 >");	// Vector No: 1492
verify(op === 'b11111111, "Assert 5969 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5970 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 5971 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111110111:0:1:1111:11111111:1:11111111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111110111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1494
#2;

verify(ir === 'b1111, "Assert 5972 : < ir !== 'b1111 >");	// Vector No: 1493
verify(op === 'b11111111, "Assert 5973 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5974 : < extop !== 1 >");
verify(addr === 'b11111111111111110111, "Assert 5975 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111110111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111110111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1495
#2;

verify(ir === 'b1111, "Assert 5976 : < ir !== 'b1111 >");	// Vector No: 1494
verify(op === 'b11111000, "Assert 5977 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5978 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5979 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111110111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111110111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1496
#2;

verify(ir === 'b1111, "Assert 5980 : < ir !== 'b1111 >");	// Vector No: 1495
verify(op === 'b11100000, "Assert 5981 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 5982 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 5983 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111110111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111110111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1497
#2;

verify(ir === 'b1111, "Assert 5984 : < ir !== 'b1111 >");	// Vector No: 1496
verify(op === 'b11111111, "Assert 5985 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 5986 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 5987 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111110111:0:1:1111:11111111:0:11111111111111110111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111110111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1498
#2;

verify(ir === 'b1111, "Assert 5988 : < ir !== 'b1111 >");	// Vector No: 1497
verify(op === 'b11111111, "Assert 5989 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 5990 : < extop !== 0 >");
verify(addr === 'b11111111111111110111, "Assert 5991 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111110111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111110111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1499
#2;

verify(ir === 'b1011, "Assert 5992 : < ir !== 'b1011 >");	// Vector No: 1498
verify(op === 'b11111000, "Assert 5993 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5994 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5995 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111110111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111110111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1500
#2;

verify(ir === 'b1111, "Assert 5996 : < ir !== 'b1111 >");	// Vector No: 1499
verify(op === 'b11111000, "Assert 5997 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 5998 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 5999 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111101111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111101111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1501
#2;

verify(ir === 'b1111, "Assert 6000 : < ir !== 'b1111 >");	// Vector No: 1500
verify(op === 'b11111111, "Assert 6001 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6002 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6003 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111101111:0:1:1111:11111111:1:11111111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111101111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1502
#2;

verify(ir === 'b1111, "Assert 6004 : < ir !== 'b1111 >");	// Vector No: 1501
verify(op === 'b11111111, "Assert 6005 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6006 : < extop !== 1 >");
verify(addr === 'b11111111111111101111, "Assert 6007 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111101111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111101111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1503
#2;

verify(ir === 'b1111, "Assert 6008 : < ir !== 'b1111 >");	// Vector No: 1502
verify(op === 'b11111000, "Assert 6009 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6010 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6011 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111101111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111101111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1504
#2;

verify(ir === 'b1111, "Assert 6012 : < ir !== 'b1111 >");	// Vector No: 1503
verify(op === 'b11100000, "Assert 6013 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6014 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6015 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111101111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111101111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1505
#2;

verify(ir === 'b1111, "Assert 6016 : < ir !== 'b1111 >");	// Vector No: 1504
verify(op === 'b11111111, "Assert 6017 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6018 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6019 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111101111:0:1:1111:11111111:0:11111111111111101111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111101111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1506
#2;

verify(ir === 'b1111, "Assert 6020 : < ir !== 'b1111 >");	// Vector No: 1505
verify(op === 'b11111111, "Assert 6021 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6022 : < extop !== 0 >");
verify(addr === 'b11111111111111101111, "Assert 6023 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111101111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111101111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1507
#2;

verify(ir === 'b1011, "Assert 6024 : < ir !== 'b1011 >");	// Vector No: 1506
verify(op === 'b11111000, "Assert 6025 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6026 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6027 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111101111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111101111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1508
#2;

verify(ir === 'b1111, "Assert 6028 : < ir !== 'b1111 >");	// Vector No: 1507
verify(op === 'b11111000, "Assert 6029 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6030 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6031 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111011111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111011111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1509
#2;

verify(ir === 'b1111, "Assert 6032 : < ir !== 'b1111 >");	// Vector No: 1508
verify(op === 'b11111111, "Assert 6033 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6034 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6035 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111011111:0:1:1111:11111111:1:11111111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111011111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1510
#2;

verify(ir === 'b1111, "Assert 6036 : < ir !== 'b1111 >");	// Vector No: 1509
verify(op === 'b11111111, "Assert 6037 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6038 : < extop !== 1 >");
verify(addr === 'b11111111111111011111, "Assert 6039 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111011111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111011111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1511
#2;

verify(ir === 'b1111, "Assert 6040 : < ir !== 'b1111 >");	// Vector No: 1510
verify(op === 'b11111000, "Assert 6041 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6042 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6043 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111011111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111011111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1512
#2;

verify(ir === 'b1111, "Assert 6044 : < ir !== 'b1111 >");	// Vector No: 1511
verify(op === 'b11100000, "Assert 6045 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6046 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6047 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111011111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111011111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1513
#2;

verify(ir === 'b1111, "Assert 6048 : < ir !== 'b1111 >");	// Vector No: 1512
verify(op === 'b11111111, "Assert 6049 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6050 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6051 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111011111:0:1:1111:11111111:0:11111111111111011111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111011111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1514
#2;

verify(ir === 'b1111, "Assert 6052 : < ir !== 'b1111 >");	// Vector No: 1513
verify(op === 'b11111111, "Assert 6053 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6054 : < extop !== 0 >");
verify(addr === 'b11111111111111011111, "Assert 6055 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111011111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111011111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1515
#2;

verify(ir === 'b1011, "Assert 6056 : < ir !== 'b1011 >");	// Vector No: 1514
verify(op === 'b11111000, "Assert 6057 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6058 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6059 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111011111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111011111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1516
#2;

verify(ir === 'b1111, "Assert 6060 : < ir !== 'b1111 >");	// Vector No: 1515
verify(op === 'b11111000, "Assert 6061 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6062 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6063 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111110111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111110111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1517
#2;

verify(ir === 'b1111, "Assert 6064 : < ir !== 'b1111 >");	// Vector No: 1516
verify(op === 'b11111111, "Assert 6065 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6066 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6067 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111110111111:0:1:1111:11111111:1:11111111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111110111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1518
#2;

verify(ir === 'b1111, "Assert 6068 : < ir !== 'b1111 >");	// Vector No: 1517
verify(op === 'b11111111, "Assert 6069 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6070 : < extop !== 1 >");
verify(addr === 'b11111111111110111111, "Assert 6071 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111110111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111110111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1519
#2;

verify(ir === 'b1111, "Assert 6072 : < ir !== 'b1111 >");	// Vector No: 1518
verify(op === 'b11111000, "Assert 6073 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6074 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6075 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111110111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111110111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1520
#2;

verify(ir === 'b1111, "Assert 6076 : < ir !== 'b1111 >");	// Vector No: 1519
verify(op === 'b11100000, "Assert 6077 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6078 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6079 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111110111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111110111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1521
#2;

verify(ir === 'b1111, "Assert 6080 : < ir !== 'b1111 >");	// Vector No: 1520
verify(op === 'b11111111, "Assert 6081 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6082 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6083 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111110111111:0:1:1111:11111111:0:11111111111110111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111110111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1522
#2;

verify(ir === 'b1111, "Assert 6084 : < ir !== 'b1111 >");	// Vector No: 1521
verify(op === 'b11111111, "Assert 6085 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6086 : < extop !== 0 >");
verify(addr === 'b11111111111110111111, "Assert 6087 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111110111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111110111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1523
#2;

verify(ir === 'b1011, "Assert 6088 : < ir !== 'b1011 >");	// Vector No: 1522
verify(op === 'b11111000, "Assert 6089 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6090 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6091 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111110111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111110111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1524
#2;

verify(ir === 'b1111, "Assert 6092 : < ir !== 'b1111 >");	// Vector No: 1523
verify(op === 'b11111000, "Assert 6093 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6094 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6095 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111101111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111101111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1525
#2;

verify(ir === 'b1111, "Assert 6096 : < ir !== 'b1111 >");	// Vector No: 1524
verify(op === 'b11111111, "Assert 6097 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6098 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6099 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111101111111:0:1:1111:11111111:1:11111111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111101111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1526
#2;

verify(ir === 'b1111, "Assert 6100 : < ir !== 'b1111 >");	// Vector No: 1525
verify(op === 'b11111111, "Assert 6101 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6102 : < extop !== 1 >");
verify(addr === 'b11111111111101111111, "Assert 6103 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111101111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111101111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1527
#2;

verify(ir === 'b1111, "Assert 6104 : < ir !== 'b1111 >");	// Vector No: 1526
verify(op === 'b11111000, "Assert 6105 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6106 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6107 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111101111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111101111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1528
#2;

verify(ir === 'b1111, "Assert 6108 : < ir !== 'b1111 >");	// Vector No: 1527
verify(op === 'b11100000, "Assert 6109 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6110 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6111 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111101111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111101111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1529
#2;

verify(ir === 'b1111, "Assert 6112 : < ir !== 'b1111 >");	// Vector No: 1528
verify(op === 'b11111111, "Assert 6113 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6114 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6115 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111101111111:0:1:1111:11111111:0:11111111111101111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111101111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1530
#2;

verify(ir === 'b1111, "Assert 6116 : < ir !== 'b1111 >");	// Vector No: 1529
verify(op === 'b11111111, "Assert 6117 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6118 : < extop !== 0 >");
verify(addr === 'b11111111111101111111, "Assert 6119 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111101111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111101111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1531
#2;

verify(ir === 'b1011, "Assert 6120 : < ir !== 'b1011 >");	// Vector No: 1530
verify(op === 'b11111000, "Assert 6121 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6122 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6123 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111101111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111101111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1532
#2;

verify(ir === 'b1111, "Assert 6124 : < ir !== 'b1111 >");	// Vector No: 1531
verify(op === 'b11111000, "Assert 6125 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6126 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6127 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111011111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111011111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1533
#2;

verify(ir === 'b1111, "Assert 6128 : < ir !== 'b1111 >");	// Vector No: 1532
verify(op === 'b11111111, "Assert 6129 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6130 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6131 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111011111111:0:1:1111:11111111:1:11111111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111011111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1534
#2;

verify(ir === 'b1111, "Assert 6132 : < ir !== 'b1111 >");	// Vector No: 1533
verify(op === 'b11111111, "Assert 6133 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6134 : < extop !== 1 >");
verify(addr === 'b11111111111011111111, "Assert 6135 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111011111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111011111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1535
#2;

verify(ir === 'b1111, "Assert 6136 : < ir !== 'b1111 >");	// Vector No: 1534
verify(op === 'b11111000, "Assert 6137 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6138 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6139 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111011111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111011111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1536
#2;

verify(ir === 'b1111, "Assert 6140 : < ir !== 'b1111 >");	// Vector No: 1535
verify(op === 'b11100000, "Assert 6141 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6142 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6143 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111011111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111011111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1537
#2;

verify(ir === 'b1111, "Assert 6144 : < ir !== 'b1111 >");	// Vector No: 1536
verify(op === 'b11111111, "Assert 6145 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6146 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6147 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111011111111:0:1:1111:11111111:0:11111111111011111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111011111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1538
#2;

verify(ir === 'b1111, "Assert 6148 : < ir !== 'b1111 >");	// Vector No: 1537
verify(op === 'b11111111, "Assert 6149 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6150 : < extop !== 0 >");
verify(addr === 'b11111111111011111111, "Assert 6151 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111011111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111011111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1539
#2;

verify(ir === 'b1011, "Assert 6152 : < ir !== 'b1011 >");	// Vector No: 1538
verify(op === 'b11111000, "Assert 6153 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6154 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6155 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111011111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111011111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1540
#2;

verify(ir === 'b1111, "Assert 6156 : < ir !== 'b1111 >");	// Vector No: 1539
verify(op === 'b11111000, "Assert 6157 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6158 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6159 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111110111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111110111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1541
#2;

verify(ir === 'b1111, "Assert 6160 : < ir !== 'b1111 >");	// Vector No: 1540
verify(op === 'b11111111, "Assert 6161 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6162 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6163 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111110111111111:0:1:1111:11111111:1:11111111110111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111110111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1542
#2;

verify(ir === 'b1111, "Assert 6164 : < ir !== 'b1111 >");	// Vector No: 1541
verify(op === 'b11111111, "Assert 6165 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6166 : < extop !== 1 >");
verify(addr === 'b11111111110111111111, "Assert 6167 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111110111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111110111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1543
#2;

verify(ir === 'b1111, "Assert 6168 : < ir !== 'b1111 >");	// Vector No: 1542
verify(op === 'b11111000, "Assert 6169 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6170 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6171 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111110111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111110111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1544
#2;

verify(ir === 'b1111, "Assert 6172 : < ir !== 'b1111 >");	// Vector No: 1543
verify(op === 'b11100000, "Assert 6173 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6174 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6175 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111110111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111110111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1545
#2;

verify(ir === 'b1111, "Assert 6176 : < ir !== 'b1111 >");	// Vector No: 1544
verify(op === 'b11111111, "Assert 6177 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6178 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6179 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111110111111111:0:1:1111:11111111:0:11111111110111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111110111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1546
#2;

verify(ir === 'b1111, "Assert 6180 : < ir !== 'b1111 >");	// Vector No: 1545
verify(op === 'b11111111, "Assert 6181 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6182 : < extop !== 0 >");
verify(addr === 'b11111111110111111111, "Assert 6183 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111110111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111110111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1547
#2;

verify(ir === 'b1011, "Assert 6184 : < ir !== 'b1011 >");	// Vector No: 1546
verify(op === 'b11111000, "Assert 6185 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6186 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6187 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111110111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111110111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1548
#2;

verify(ir === 'b1111, "Assert 6188 : < ir !== 'b1111 >");	// Vector No: 1547
verify(op === 'b11111000, "Assert 6189 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6190 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6191 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111101111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111101111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1549
#2;

verify(ir === 'b1111, "Assert 6192 : < ir !== 'b1111 >");	// Vector No: 1548
verify(op === 'b11111111, "Assert 6193 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6194 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6195 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111101111111111:0:1:1111:11111111:1:11111111101111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111101111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1550
#2;

verify(ir === 'b1111, "Assert 6196 : < ir !== 'b1111 >");	// Vector No: 1549
verify(op === 'b11111111, "Assert 6197 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6198 : < extop !== 1 >");
verify(addr === 'b11111111101111111111, "Assert 6199 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111101111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111101111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1551
#2;

verify(ir === 'b1111, "Assert 6200 : < ir !== 'b1111 >");	// Vector No: 1550
verify(op === 'b11111000, "Assert 6201 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6202 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6203 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111101111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111101111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1552
#2;

verify(ir === 'b1111, "Assert 6204 : < ir !== 'b1111 >");	// Vector No: 1551
verify(op === 'b11100000, "Assert 6205 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6206 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6207 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111101111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111101111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1553
#2;

verify(ir === 'b1111, "Assert 6208 : < ir !== 'b1111 >");	// Vector No: 1552
verify(op === 'b11111111, "Assert 6209 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6210 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6211 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111101111111111:0:1:1111:11111111:0:11111111101111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111101111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1554
#2;

verify(ir === 'b1111, "Assert 6212 : < ir !== 'b1111 >");	// Vector No: 1553
verify(op === 'b11111111, "Assert 6213 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6214 : < extop !== 0 >");
verify(addr === 'b11111111101111111111, "Assert 6215 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111101111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111101111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1555
#2;

verify(ir === 'b1011, "Assert 6216 : < ir !== 'b1011 >");	// Vector No: 1554
verify(op === 'b11111000, "Assert 6217 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6218 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6219 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111101111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111101111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1556
#2;

verify(ir === 'b1111, "Assert 6220 : < ir !== 'b1111 >");	// Vector No: 1555
verify(op === 'b11111000, "Assert 6221 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6222 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6223 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111011111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111011111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1557
#2;

verify(ir === 'b1111, "Assert 6224 : < ir !== 'b1111 >");	// Vector No: 1556
verify(op === 'b11111111, "Assert 6225 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6226 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6227 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111011111111111:0:1:1111:11111111:1:11111111011111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111011111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1558
#2;

verify(ir === 'b1111, "Assert 6228 : < ir !== 'b1111 >");	// Vector No: 1557
verify(op === 'b11111111, "Assert 6229 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6230 : < extop !== 1 >");
verify(addr === 'b11111111011111111111, "Assert 6231 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111011111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111011111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1559
#2;

verify(ir === 'b1111, "Assert 6232 : < ir !== 'b1111 >");	// Vector No: 1558
verify(op === 'b11111000, "Assert 6233 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6234 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6235 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111011111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111011111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1560
#2;

verify(ir === 'b1111, "Assert 6236 : < ir !== 'b1111 >");	// Vector No: 1559
verify(op === 'b11100000, "Assert 6237 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6238 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6239 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111011111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111011111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1561
#2;

verify(ir === 'b1111, "Assert 6240 : < ir !== 'b1111 >");	// Vector No: 1560
verify(op === 'b11111111, "Assert 6241 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6242 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6243 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111011111111111:0:1:1111:11111111:0:11111111011111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111011111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1562
#2;

verify(ir === 'b1111, "Assert 6244 : < ir !== 'b1111 >");	// Vector No: 1561
verify(op === 'b11111111, "Assert 6245 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6246 : < extop !== 0 >");
verify(addr === 'b11111111011111111111, "Assert 6247 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111011111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111011111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1563
#2;

verify(ir === 'b1011, "Assert 6248 : < ir !== 'b1011 >");	// Vector No: 1562
verify(op === 'b11111000, "Assert 6249 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6250 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6251 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111011111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111011111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1564
#2;

verify(ir === 'b1111, "Assert 6252 : < ir !== 'b1111 >");	// Vector No: 1563
verify(op === 'b11111000, "Assert 6253 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6254 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6255 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111110111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111110111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1565
#2;

verify(ir === 'b1111, "Assert 6256 : < ir !== 'b1111 >");	// Vector No: 1564
verify(op === 'b11111111, "Assert 6257 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6258 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6259 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111110111111111111:0:1:1111:11111110:1:11111110111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111110111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1566
#2;

verify(ir === 'b1111, "Assert 6260 : < ir !== 'b1111 >");	// Vector No: 1565
verify(op === 'b11111110, "Assert 6261 : < op !== 'b11111110 >");
verify(extop === 1, "Assert 6262 : < extop !== 1 >");
verify(addr === 'b11111110111111111111, "Assert 6263 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111110111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111110111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1567
#2;

verify(ir === 'b1111, "Assert 6264 : < ir !== 'b1111 >");	// Vector No: 1566
verify(op === 'b11111000, "Assert 6265 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6266 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6267 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111110111111111111:1:1:1111:11100000:0:00000011111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111110111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1568
#2;

verify(ir === 'b1111, "Assert 6268 : < ir !== 'b1111 >");	// Vector No: 1567
verify(op === 'b11100000, "Assert 6269 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6270 : < extop !== 0 >");
verify(addr === 'b00000011111111111110, "Assert 6271 : < addr !== 'b00000011111111111110 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111110111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111110111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1569
#2;

verify(ir === 'b1111, "Assert 6272 : < ir !== 'b1111 >");	// Vector No: 1568
verify(op === 'b11111111, "Assert 6273 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6274 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6275 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111110111111111111:0:1:1111:11111111:0:11111110111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111110111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1570
#2;

verify(ir === 'b1111, "Assert 6276 : < ir !== 'b1111 >");	// Vector No: 1569
verify(op === 'b11111111, "Assert 6277 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6278 : < extop !== 0 >");
verify(addr === 'b11111110111111111111, "Assert 6279 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111110111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111110111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1571
#2;

verify(ir === 'b1011, "Assert 6280 : < ir !== 'b1011 >");	// Vector No: 1570
verify(op === 'b11111000, "Assert 6281 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6282 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6283 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111110111111111111:1:1:1111:11111000:0:00000111111111111110:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111110111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1572
#2;

verify(ir === 'b1111, "Assert 6284 : < ir !== 'b1111 >");	// Vector No: 1571
verify(op === 'b11111000, "Assert 6285 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6286 : < extop !== 0 >");
verify(addr === 'b00000111111111111110, "Assert 6287 : < addr !== 'b00000111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111101111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111101111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1573
#2;

verify(ir === 'b1111, "Assert 6288 : < ir !== 'b1111 >");	// Vector No: 1572
verify(op === 'b11111111, "Assert 6289 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6290 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6291 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111101111111111111:0:1:1111:11111101:1:11111101111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111101111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1574
#2;

verify(ir === 'b1111, "Assert 6292 : < ir !== 'b1111 >");	// Vector No: 1573
verify(op === 'b11111101, "Assert 6293 : < op !== 'b11111101 >");
verify(extop === 1, "Assert 6294 : < extop !== 1 >");
verify(addr === 'b11111101111111111111, "Assert 6295 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111101111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111101111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1575
#2;

verify(ir === 'b1111, "Assert 6296 : < ir !== 'b1111 >");	// Vector No: 1574
verify(op === 'b11111000, "Assert 6297 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6298 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6299 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111101111111111111:1:1:1111:11100000:0:00000011111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111101111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1576
#2;

verify(ir === 'b1111, "Assert 6300 : < ir !== 'b1111 >");	// Vector No: 1575
verify(op === 'b11100000, "Assert 6301 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6302 : < extop !== 0 >");
verify(addr === 'b00000011111111111101, "Assert 6303 : < addr !== 'b00000011111111111101 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111101111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111101111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1577
#2;

verify(ir === 'b1111, "Assert 6304 : < ir !== 'b1111 >");	// Vector No: 1576
verify(op === 'b11111111, "Assert 6305 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6306 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6307 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111101111111111111:0:1:1111:11111111:0:11111101111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111101111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1578
#2;

verify(ir === 'b1111, "Assert 6308 : < ir !== 'b1111 >");	// Vector No: 1577
verify(op === 'b11111111, "Assert 6309 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6310 : < extop !== 0 >");
verify(addr === 'b11111101111111111111, "Assert 6311 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111101111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111101111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1579
#2;

verify(ir === 'b1011, "Assert 6312 : < ir !== 'b1011 >");	// Vector No: 1578
verify(op === 'b11111000, "Assert 6313 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6314 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6315 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111101111111111111:1:1:1111:11111000:0:00000111111111111101:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111101111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1580
#2;

verify(ir === 'b1111, "Assert 6316 : < ir !== 'b1111 >");	// Vector No: 1579
verify(op === 'b11111000, "Assert 6317 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6318 : < extop !== 0 >");
verify(addr === 'b00000111111111111101, "Assert 6319 : < addr !== 'b00000111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111011111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111011111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1581
#2;

verify(ir === 'b1111, "Assert 6320 : < ir !== 'b1111 >");	// Vector No: 1580
verify(op === 'b11111111, "Assert 6321 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6322 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6323 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111011111111111111:0:1:1111:11111011:1:11111011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111011111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1582
#2;

verify(ir === 'b1111, "Assert 6324 : < ir !== 'b1111 >");	// Vector No: 1581
verify(op === 'b11111011, "Assert 6325 : < op !== 'b11111011 >");
verify(extop === 1, "Assert 6326 : < extop !== 1 >");
verify(addr === 'b11111011111111111111, "Assert 6327 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111011111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111011111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1583
#2;

verify(ir === 'b1111, "Assert 6328 : < ir !== 'b1111 >");	// Vector No: 1582
verify(op === 'b11111000, "Assert 6329 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6330 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6331 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111011111111111111:1:1:1111:11100000:0:00000011111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111011111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1584
#2;

verify(ir === 'b1111, "Assert 6332 : < ir !== 'b1111 >");	// Vector No: 1583
verify(op === 'b11100000, "Assert 6333 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6334 : < extop !== 0 >");
verify(addr === 'b00000011111111111011, "Assert 6335 : < addr !== 'b00000011111111111011 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111011111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111011111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1585
#2;

verify(ir === 'b1111, "Assert 6336 : < ir !== 'b1111 >");	// Vector No: 1584
verify(op === 'b11111111, "Assert 6337 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6338 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6339 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111011111111111111:0:1:1111:11111111:0:11111011111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111011111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1586
#2;

verify(ir === 'b1111, "Assert 6340 : < ir !== 'b1111 >");	// Vector No: 1585
verify(op === 'b11111111, "Assert 6341 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6342 : < extop !== 0 >");
verify(addr === 'b11111011111111111111, "Assert 6343 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111011111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111011111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1587
#2;

verify(ir === 'b1011, "Assert 6344 : < ir !== 'b1011 >");	// Vector No: 1586
verify(op === 'b11111000, "Assert 6345 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6346 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6347 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111011111111111111:1:1:1111:11111000:0:00000111111111111011:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111011111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1588
#2;

verify(ir === 'b1111, "Assert 6348 : < ir !== 'b1111 >");	// Vector No: 1587
verify(op === 'b11111000, "Assert 6349 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6350 : < extop !== 0 >");
verify(addr === 'b00000111111111111011, "Assert 6351 : < addr !== 'b00000111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111110111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111110111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1589
#2;

verify(ir === 'b1111, "Assert 6352 : < ir !== 'b1111 >");	// Vector No: 1588
verify(op === 'b11111111, "Assert 6353 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6354 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6355 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111110111111111111111:0:1:1111:11110111:1:11110111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111110111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1590
#2;

verify(ir === 'b1111, "Assert 6356 : < ir !== 'b1111 >");	// Vector No: 1589
verify(op === 'b11110111, "Assert 6357 : < op !== 'b11110111 >");
verify(extop === 1, "Assert 6358 : < extop !== 1 >");
verify(addr === 'b11110111111111111111, "Assert 6359 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111110111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111110111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1591
#2;

verify(ir === 'b1111, "Assert 6360 : < ir !== 'b1111 >");	// Vector No: 1590
verify(op === 'b11111000, "Assert 6361 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6362 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6363 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111110111111111111111:1:1:1111:11100000:0:00000011111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111110111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1592
#2;

verify(ir === 'b1111, "Assert 6364 : < ir !== 'b1111 >");	// Vector No: 1591
verify(op === 'b11100000, "Assert 6365 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6366 : < extop !== 0 >");
verify(addr === 'b00000011111111110111, "Assert 6367 : < addr !== 'b00000011111111110111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111110111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111110111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1593
#2;

verify(ir === 'b1111, "Assert 6368 : < ir !== 'b1111 >");	// Vector No: 1592
verify(op === 'b11111111, "Assert 6369 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6370 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6371 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111110111111111111111:0:1:1111:11111111:0:11110111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111110111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1594
#2;

verify(ir === 'b1111, "Assert 6372 : < ir !== 'b1111 >");	// Vector No: 1593
verify(op === 'b11111111, "Assert 6373 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6374 : < extop !== 0 >");
verify(addr === 'b11110111111111111111, "Assert 6375 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111110111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111110111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1595
#2;

verify(ir === 'b1011, "Assert 6376 : < ir !== 'b1011 >");	// Vector No: 1594
verify(op === 'b11111000, "Assert 6377 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6378 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6379 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111110111111111111111:1:1:1111:11111000:0:00000111111111110111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111110111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1596
#2;

verify(ir === 'b1111, "Assert 6380 : < ir !== 'b1111 >");	// Vector No: 1595
verify(op === 'b11111000, "Assert 6381 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6382 : < extop !== 0 >");
verify(addr === 'b00000111111111110111, "Assert 6383 : < addr !== 'b00000111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111101111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111101111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1597
#2;

verify(ir === 'b1111, "Assert 6384 : < ir !== 'b1111 >");	// Vector No: 1596
verify(op === 'b11111111, "Assert 6385 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6386 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6387 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111101111111111111111:0:1:1111:11101111:1:11101111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111101111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1598
#2;

verify(ir === 'b1111, "Assert 6388 : < ir !== 'b1111 >");	// Vector No: 1597
verify(op === 'b11101111, "Assert 6389 : < op !== 'b11101111 >");
verify(extop === 1, "Assert 6390 : < extop !== 1 >");
verify(addr === 'b11101111111111111111, "Assert 6391 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111101111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111101111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1599
#2;

verify(ir === 'b1111, "Assert 6392 : < ir !== 'b1111 >");	// Vector No: 1598
verify(op === 'b11111000, "Assert 6393 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6394 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6395 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111101111111111111111:1:1:1111:11100000:0:00000011111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111101111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1600
#2;

verify(ir === 'b1111, "Assert 6396 : < ir !== 'b1111 >");	// Vector No: 1599
verify(op === 'b11100000, "Assert 6397 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6398 : < extop !== 0 >");
verify(addr === 'b00000011111111101111, "Assert 6399 : < addr !== 'b00000011111111101111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111101111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111101111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1601
#2;

verify(ir === 'b1111, "Assert 6400 : < ir !== 'b1111 >");	// Vector No: 1600
verify(op === 'b11111111, "Assert 6401 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6402 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6403 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111101111111111111111:0:1:1111:11111111:0:11101111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111101111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1602
#2;

verify(ir === 'b1111, "Assert 6404 : < ir !== 'b1111 >");	// Vector No: 1601
verify(op === 'b11111111, "Assert 6405 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6406 : < extop !== 0 >");
verify(addr === 'b11101111111111111111, "Assert 6407 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111101111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111101111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1603
#2;

verify(ir === 'b1011, "Assert 6408 : < ir !== 'b1011 >");	// Vector No: 1602
verify(op === 'b11111000, "Assert 6409 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6410 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6411 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111101111111111111111:1:1:1111:11111000:0:00000111111111101111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111101111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1604
#2;

verify(ir === 'b1111, "Assert 6412 : < ir !== 'b1111 >");	// Vector No: 1603
verify(op === 'b11111000, "Assert 6413 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6414 : < extop !== 0 >");
verify(addr === 'b00000111111111101111, "Assert 6415 : < addr !== 'b00000111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111011111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111011111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1605
#2;

verify(ir === 'b1111, "Assert 6416 : < ir !== 'b1111 >");	// Vector No: 1604
verify(op === 'b11111111, "Assert 6417 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6418 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6419 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111011111111111111111:0:1:1111:11011111:1:11011111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111011111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1606
#2;

verify(ir === 'b1111, "Assert 6420 : < ir !== 'b1111 >");	// Vector No: 1605
verify(op === 'b11011111, "Assert 6421 : < op !== 'b11011111 >");
verify(extop === 1, "Assert 6422 : < extop !== 1 >");
verify(addr === 'b11011111111111111111, "Assert 6423 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111011111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111011111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1607
#2;

verify(ir === 'b1111, "Assert 6424 : < ir !== 'b1111 >");	// Vector No: 1606
verify(op === 'b11111000, "Assert 6425 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6426 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6427 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111011111111111111111:1:1:1111:11100000:0:00000011111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111011111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1608
#2;

verify(ir === 'b1111, "Assert 6428 : < ir !== 'b1111 >");	// Vector No: 1607
verify(op === 'b11100000, "Assert 6429 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6430 : < extop !== 0 >");
verify(addr === 'b00000011111111011111, "Assert 6431 : < addr !== 'b00000011111111011111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111011111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111011111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1609
#2;

verify(ir === 'b1111, "Assert 6432 : < ir !== 'b1111 >");	// Vector No: 1608
verify(op === 'b11111111, "Assert 6433 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6434 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6435 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111011111111111111111:0:1:1111:11111111:0:11011111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111011111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1610
#2;

verify(ir === 'b1111, "Assert 6436 : < ir !== 'b1111 >");	// Vector No: 1609
verify(op === 'b11111111, "Assert 6437 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6438 : < extop !== 0 >");
verify(addr === 'b11011111111111111111, "Assert 6439 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111011111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111011111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1611
#2;

verify(ir === 'b1011, "Assert 6440 : < ir !== 'b1011 >");	// Vector No: 1610
verify(op === 'b11111000, "Assert 6441 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6442 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6443 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111011111111111111111:1:1:1111:11111000:0:00000111111111011111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111011111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1612
#2;

verify(ir === 'b1111, "Assert 6444 : < ir !== 'b1111 >");	// Vector No: 1611
verify(op === 'b11111000, "Assert 6445 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6446 : < extop !== 0 >");
verify(addr === 'b00000111111111011111, "Assert 6447 : < addr !== 'b00000111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111110111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111110111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1613
#2;

verify(ir === 'b1111, "Assert 6448 : < ir !== 'b1111 >");	// Vector No: 1612
verify(op === 'b11111111, "Assert 6449 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6450 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6451 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111110111111111111111111:0:1:1111:10111111:1:10111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111110111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1614
#2;

verify(ir === 'b1111, "Assert 6452 : < ir !== 'b1111 >");	// Vector No: 1613
verify(op === 'b10111111, "Assert 6453 : < op !== 'b10111111 >");
verify(extop === 1, "Assert 6454 : < extop !== 1 >");
verify(addr === 'b10111111111111111111, "Assert 6455 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111110111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111110111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1615
#2;

verify(ir === 'b1111, "Assert 6456 : < ir !== 'b1111 >");	// Vector No: 1614
verify(op === 'b11111000, "Assert 6457 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6458 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6459 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111110111111111111111111:1:1:1111:11100000:0:00000011111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111110111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1616
#2;

verify(ir === 'b1111, "Assert 6460 : < ir !== 'b1111 >");	// Vector No: 1615
verify(op === 'b11100000, "Assert 6461 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6462 : < extop !== 0 >");
verify(addr === 'b00000011111110111111, "Assert 6463 : < addr !== 'b00000011111110111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111110111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111110111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1617
#2;

verify(ir === 'b1111, "Assert 6464 : < ir !== 'b1111 >");	// Vector No: 1616
verify(op === 'b11111111, "Assert 6465 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6466 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6467 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111110111111111111111111:0:1:1111:11111111:0:10111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111110111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1618
#2;

verify(ir === 'b1111, "Assert 6468 : < ir !== 'b1111 >");	// Vector No: 1617
verify(op === 'b11111111, "Assert 6469 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6470 : < extop !== 0 >");
verify(addr === 'b10111111111111111111, "Assert 6471 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111110111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111110111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1619
#2;

verify(ir === 'b1011, "Assert 6472 : < ir !== 'b1011 >");	// Vector No: 1618
verify(op === 'b11111000, "Assert 6473 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6474 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6475 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111110111111111111111111:1:1:1111:11111000:0:00000111111110111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111110111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1620
#2;

verify(ir === 'b1111, "Assert 6476 : < ir !== 'b1111 >");	// Vector No: 1619
verify(op === 'b11111000, "Assert 6477 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6478 : < extop !== 0 >");
verify(addr === 'b00000111111110111111, "Assert 6479 : < addr !== 'b00000111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111101111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111101111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1621
#2;

verify(ir === 'b1111, "Assert 6480 : < ir !== 'b1111 >");	// Vector No: 1620
verify(op === 'b11111111, "Assert 6481 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6482 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6483 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111101111111111111111111:0:1:1111:01111111:1:01111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111101111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1622
#2;

verify(ir === 'b1111, "Assert 6484 : < ir !== 'b1111 >");	// Vector No: 1621
verify(op === 'b01111111, "Assert 6485 : < op !== 'b01111111 >");
verify(extop === 1, "Assert 6486 : < extop !== 1 >");
verify(addr === 'b01111111111111111111, "Assert 6487 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111101111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111101111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1623
#2;

verify(ir === 'b1111, "Assert 6488 : < ir !== 'b1111 >");	// Vector No: 1622
verify(op === 'b11111000, "Assert 6489 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6490 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6491 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111101111111111111111111:1:1:1111:11100000:0:00000011111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111101111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1624
#2;

verify(ir === 'b1111, "Assert 6492 : < ir !== 'b1111 >");	// Vector No: 1623
verify(op === 'b11100000, "Assert 6493 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6494 : < extop !== 0 >");
verify(addr === 'b00000011111101111111, "Assert 6495 : < addr !== 'b00000011111101111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111101111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111101111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1625
#2;

verify(ir === 'b1111, "Assert 6496 : < ir !== 'b1111 >");	// Vector No: 1624
verify(op === 'b11111111, "Assert 6497 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6498 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6499 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111101111111111111111111:0:1:1111:11111111:0:01111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111101111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1626
#2;

verify(ir === 'b1111, "Assert 6500 : < ir !== 'b1111 >");	// Vector No: 1625
verify(op === 'b11111111, "Assert 6501 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6502 : < extop !== 0 >");
verify(addr === 'b01111111111111111111, "Assert 6503 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111101111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111101111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1627
#2;

verify(ir === 'b1011, "Assert 6504 : < ir !== 'b1011 >");	// Vector No: 1626
verify(op === 'b11111000, "Assert 6505 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6506 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6507 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111101111111111111111111:1:1:1111:11111000:0:00000111111101111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111101111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1628
#2;

verify(ir === 'b1111, "Assert 6508 : < ir !== 'b1111 >");	// Vector No: 1627
verify(op === 'b11111000, "Assert 6509 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6510 : < extop !== 0 >");
verify(addr === 'b00000111111101111111, "Assert 6511 : < addr !== 'b00000111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1629
#2;

verify(ir === 'b1111, "Assert 6512 : < ir !== 'b1111 >");	// Vector No: 1628
verify(op === 'b11111111, "Assert 6513 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6514 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6515 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1630
#2;

verify(ir === 'b1111, "Assert 6516 : < ir !== 'b1111 >");	// Vector No: 1629
verify(op === 'b11111111, "Assert 6517 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6518 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6519 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1631
#2;

verify(ir === 'b1111, "Assert 6520 : < ir !== 'b1111 >");	// Vector No: 1630
verify(op === 'b11111000, "Assert 6521 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6522 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6523 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1632
#2;

verify(ir === 'b1111, "Assert 6524 : < ir !== 'b1111 >");	// Vector No: 1631
verify(op === 'b11100000, "Assert 6525 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6526 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6527 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111011111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111011111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1633
#2;

verify(ir === 'b1111, "Assert 6528 : < ir !== 'b1111 >");	// Vector No: 1632
verify(op === 'b11111111, "Assert 6529 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6530 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6531 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111011111111111111111111:0:1:1111:11111110:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111011111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1634
#2;

verify(ir === 'b1111, "Assert 6532 : < ir !== 'b1111 >");	// Vector No: 1633
verify(op === 'b11111110, "Assert 6533 : < op !== 'b11111110 >");
verify(extop === 0, "Assert 6534 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6535 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111011111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111011111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1635
#2;

verify(ir === 'b1011, "Assert 6536 : < ir !== 'b1011 >");	// Vector No: 1634
verify(op === 'b11111000, "Assert 6537 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6538 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6539 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111011111111111111111111:1:1:1111:11111000:0:00000111111011111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111011111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1636
#2;

verify(ir === 'b1111, "Assert 6540 : < ir !== 'b1111 >");	// Vector No: 1635
verify(op === 'b11111000, "Assert 6541 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6542 : < extop !== 0 >");
verify(addr === 'b00000111111011111111, "Assert 6543 : < addr !== 'b00000111111011111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111110111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111110111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1637
#2;

verify(ir === 'b1111, "Assert 6544 : < ir !== 'b1111 >");	// Vector No: 1636
verify(op === 'b11111111, "Assert 6545 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6546 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6547 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111110111111111111111111111:0:1:1111:11111101:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111110111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1638
#2;

verify(ir === 'b1111, "Assert 6548 : < ir !== 'b1111 >");	// Vector No: 1637
verify(op === 'b11111101, "Assert 6549 : < op !== 'b11111101 >");
verify(extop === 0, "Assert 6550 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6551 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111110111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111110111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1639
#2;

verify(ir === 'b1011, "Assert 6552 : < ir !== 'b1011 >");	// Vector No: 1638
verify(op === 'b11111000, "Assert 6553 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6554 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6555 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111110111111111111111111111:1:1:1111:11111000:0:00000111110111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111110111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1640
#2;

verify(ir === 'b1111, "Assert 6556 : < ir !== 'b1111 >");	// Vector No: 1639
verify(op === 'b11111000, "Assert 6557 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6558 : < extop !== 0 >");
verify(addr === 'b00000111110111111111, "Assert 6559 : < addr !== 'b00000111110111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111101111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111101111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1641
#2;

verify(ir === 'b1111, "Assert 6560 : < ir !== 'b1111 >");	// Vector No: 1640
verify(op === 'b11111111, "Assert 6561 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6562 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6563 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111101111111111111111111111:0:1:1111:11111011:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111101111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1642
#2;

verify(ir === 'b1111, "Assert 6564 : < ir !== 'b1111 >");	// Vector No: 1641
verify(op === 'b11111011, "Assert 6565 : < op !== 'b11111011 >");
verify(extop === 0, "Assert 6566 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6567 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111101111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111101111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1643
#2;

verify(ir === 'b1011, "Assert 6568 : < ir !== 'b1011 >");	// Vector No: 1642
verify(op === 'b11111000, "Assert 6569 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6570 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6571 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111101111111111111111111111:1:1:1111:11111000:0:00000111101111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111101111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1644
#2;

verify(ir === 'b1111, "Assert 6572 : < ir !== 'b1111 >");	// Vector No: 1643
verify(op === 'b11111000, "Assert 6573 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6574 : < extop !== 0 >");
verify(addr === 'b00000111101111111111, "Assert 6575 : < addr !== 'b00000111101111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111011111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111011111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1645
#2;

verify(ir === 'b1111, "Assert 6576 : < ir !== 'b1111 >");	// Vector No: 1644
verify(op === 'b11111111, "Assert 6577 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6578 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6579 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111011111111111111111111111:0:1:1111:11110111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111011111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1646
#2;

verify(ir === 'b1111, "Assert 6580 : < ir !== 'b1111 >");	// Vector No: 1645
verify(op === 'b11110111, "Assert 6581 : < op !== 'b11110111 >");
verify(extop === 0, "Assert 6582 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6583 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111011111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111011111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1647
#2;

verify(ir === 'b1011, "Assert 6584 : < ir !== 'b1011 >");	// Vector No: 1646
verify(op === 'b11111000, "Assert 6585 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6586 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6587 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111011111111111111111111111:1:1:1111:11111000:0:00000111011111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111011111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1648
#2;

verify(ir === 'b1111, "Assert 6588 : < ir !== 'b1111 >");	// Vector No: 1647
verify(op === 'b11111000, "Assert 6589 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6590 : < extop !== 0 >");
verify(addr === 'b00000111011111111111, "Assert 6591 : < addr !== 'b00000111011111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111110111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111110111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1649
#2;

verify(ir === 'b1111, "Assert 6592 : < ir !== 'b1111 >");	// Vector No: 1648
verify(op === 'b11111111, "Assert 6593 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6594 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6595 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111110111111111111111111111111:0:1:1111:11101111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111110111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1650
#2;

verify(ir === 'b1111, "Assert 6596 : < ir !== 'b1111 >");	// Vector No: 1649
verify(op === 'b11101111, "Assert 6597 : < op !== 'b11101111 >");
verify(extop === 0, "Assert 6598 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6599 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111110111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111110111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1651
#2;

verify(ir === 'b1011, "Assert 6600 : < ir !== 'b1011 >");	// Vector No: 1650
verify(op === 'b11111000, "Assert 6601 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6602 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6603 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111110111111111111111111111111:1:1:1111:11111000:0:00000110111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111110111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1652
#2;

verify(ir === 'b1111, "Assert 6604 : < ir !== 'b1111 >");	// Vector No: 1651
verify(op === 'b11111000, "Assert 6605 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6606 : < extop !== 0 >");
verify(addr === 'b00000110111111111111, "Assert 6607 : < addr !== 'b00000110111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111101111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111101111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1653
#2;

verify(ir === 'b1111, "Assert 6608 : < ir !== 'b1111 >");	// Vector No: 1652
verify(op === 'b11111111, "Assert 6609 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6610 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6611 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111101111111111111111111111111:0:1:1111:11011111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111101111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1654
#2;

verify(ir === 'b1111, "Assert 6612 : < ir !== 'b1111 >");	// Vector No: 1653
verify(op === 'b11011111, "Assert 6613 : < op !== 'b11011111 >");
verify(extop === 0, "Assert 6614 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6615 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111101111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111101111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1655
#2;

verify(ir === 'b1011, "Assert 6616 : < ir !== 'b1011 >");	// Vector No: 1654
verify(op === 'b11111000, "Assert 6617 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6618 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6619 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111101111111111111111111111111:1:1:1111:11111000:0:00000101111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111101111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1656
#2;

verify(ir === 'b1111, "Assert 6620 : < ir !== 'b1111 >");	// Vector No: 1655
verify(op === 'b11111000, "Assert 6621 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6622 : < extop !== 0 >");
verify(addr === 'b00000101111111111111, "Assert 6623 : < addr !== 'b00000101111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111011111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1657
#2;

verify(ir === 'b1111, "Assert 6624 : < ir !== 'b1111 >");	// Vector No: 1656
verify(op === 'b11111111, "Assert 6625 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6626 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6627 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111011111111111111111111111111:0:1:1111:10111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1658
#2;

verify(ir === 'b1111, "Assert 6628 : < ir !== 'b1111 >");	// Vector No: 1657
verify(op === 'b10111111, "Assert 6629 : < op !== 'b10111111 >");
verify(extop === 0, "Assert 6630 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6631 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111011111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1659
#2;

verify(ir === 'b1011, "Assert 6632 : < ir !== 'b1011 >");	// Vector No: 1658
verify(op === 'b11111000, "Assert 6633 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6634 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6635 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111011111111111111111111111111:1:1:1111:11110000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1660
#2;

verify(ir === 'b1111, "Assert 6636 : < ir !== 'b1111 >");	// Vector No: 1659
verify(op === 'b11110000, "Assert 6637 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 6638 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6639 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111110111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111110111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1661
#2;

verify(ir === 'b1111, "Assert 6640 : < ir !== 'b1111 >");	// Vector No: 1660
verify(op === 'b11111111, "Assert 6641 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6642 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6643 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111110111111111111111111111111111:0:1:1111:01111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111110111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1662
#2;

verify(ir === 'b1111, "Assert 6644 : < ir !== 'b1111 >");	// Vector No: 1661
verify(op === 'b01111111, "Assert 6645 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 6646 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6647 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111110111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111110111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1663
#2;

verify(ir === 'b1011, "Assert 6648 : < ir !== 'b1011 >");	// Vector No: 1662
verify(op === 'b11111000, "Assert 6649 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6650 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6651 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111110111111111111111111111111111:1:1:1111:11101000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111110111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1664
#2;

verify(ir === 'b1111, "Assert 6652 : < ir !== 'b1111 >");	// Vector No: 1663
verify(op === 'b11101000, "Assert 6653 : < op !== 'b11101000 >");
verify(extop === 0, "Assert 6654 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6655 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111100011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111100011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1665
#2;

verify(ir === 'b1111, "Assert 6656 : < ir !== 'b1111 >");	// Vector No: 1664
verify(op === 'b11111111, "Assert 6657 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6658 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6659 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111100011111111111111111111111111:0:1:1110:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111100011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1666
#2;

verify(ir === 'b1110, "Assert 6660 : < ir !== 'b1110 >");	// Vector No: 1665
verify(op === 'b11111111, "Assert 6661 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6662 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6663 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111100011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111100011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1667
#2;

verify(ir === 'b1111, "Assert 6664 : < ir !== 'b1111 >");	// Vector No: 1666
verify(op === 'b11111000, "Assert 6665 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6666 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6667 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111100011111111111111111111111111:1:1:1111:11000000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111100011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1668
#2;

verify(ir === 'b1111, "Assert 6668 : < ir !== 'b1111 >");	// Vector No: 1667
verify(op === 'b11000000, "Assert 6669 : < op !== 'b11000000 >");
verify(extop === 0, "Assert 6670 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6671 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111101111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111101111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1669
#2;

verify(ir === 'b1111, "Assert 6672 : < ir !== 'b1111 >");	// Vector No: 1668
verify(op === 'b11111111, "Assert 6673 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6674 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6675 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111101111111111111111111111111111:0:1:1110:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111101111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1670
#2;

verify(ir === 'b1110, "Assert 6676 : < ir !== 'b1110 >");	// Vector No: 1669
verify(op === 'b11111111, "Assert 6677 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6678 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6679 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111101111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111101111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1671
#2;

verify(ir === 'b1011, "Assert 6680 : < ir !== 'b1011 >");	// Vector No: 1670
verify(op === 'b11111000, "Assert 6681 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6682 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6683 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111101111111111111111111111111111:1:1:1111:11011000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111101111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1672
#2;

verify(ir === 'b1111, "Assert 6684 : < ir !== 'b1111 >");	// Vector No: 1671
verify(op === 'b11011000, "Assert 6685 : < op !== 'b11011000 >");
verify(extop === 0, "Assert 6686 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6687 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111010011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111010011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1673
#2;

verify(ir === 'b1111, "Assert 6688 : < ir !== 'b1111 >");	// Vector No: 1672
verify(op === 'b11111111, "Assert 6689 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6690 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6691 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111010011111111111111111111111111:0:1:1101:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111010011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1674
#2;

verify(ir === 'b1101, "Assert 6692 : < ir !== 'b1101 >");	// Vector No: 1673
verify(op === 'b11111111, "Assert 6693 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6694 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6695 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111010011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111010011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1675
#2;

verify(ir === 'b1111, "Assert 6696 : < ir !== 'b1111 >");	// Vector No: 1674
verify(op === 'b11111000, "Assert 6697 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6698 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6699 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111111010011111111111111111111111111:1:1:1111:10100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111111010011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1676
#2;

verify(ir === 'b1111, "Assert 6700 : < ir !== 'b1111 >");	// Vector No: 1675
verify(op === 'b10100000, "Assert 6701 : < op !== 'b10100000 >");
verify(extop === 0, "Assert 6702 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6703 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111011111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111011111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1677
#2;

verify(ir === 'b1111, "Assert 6704 : < ir !== 'b1111 >");	// Vector No: 1676
verify(op === 'b11111111, "Assert 6705 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6706 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6707 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111011111111111111111111111111111:0:1:1101:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111011111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1678
#2;

verify(ir === 'b1101, "Assert 6708 : < ir !== 'b1101 >");	// Vector No: 1677
verify(op === 'b11111111, "Assert 6709 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6710 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6711 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111011111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111011111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1679
#2;

verify(ir === 'b1011, "Assert 6712 : < ir !== 'b1011 >");	// Vector No: 1678
verify(op === 'b11111000, "Assert 6713 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6714 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6715 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111011111111111111111111111111111:1:1:1111:10111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111011111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1680
#2;

verify(ir === 'b1111, "Assert 6716 : < ir !== 'b1111 >");	// Vector No: 1679
verify(op === 'b10111000, "Assert 6717 : < op !== 'b10111000 >");
verify(extop === 0, "Assert 6718 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6719 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1681
#2;

verify(ir === 'b1111, "Assert 6720 : < ir !== 'b1111 >");	// Vector No: 1680
verify(op === 'b11111111, "Assert 6721 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6722 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6723 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110110011111111111111111111111111:0:1:1011:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1682
#2;

verify(ir === 'b1011, "Assert 6724 : < ir !== 'b1011 >");	// Vector No: 1681
verify(op === 'b11111111, "Assert 6725 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6726 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6727 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1683
#2;

verify(ir === 'b1111, "Assert 6728 : < ir !== 'b1111 >");	// Vector No: 1682
verify(op === 'b11111000, "Assert 6729 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6730 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6731 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111110110011111111111111111111111111:1:1:1111:01100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111110110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1684
#2;

verify(ir === 'b1111, "Assert 6732 : < ir !== 'b1111 >");	// Vector No: 1683
verify(op === 'b01100000, "Assert 6733 : < op !== 'b01100000 >");
verify(extop === 0, "Assert 6734 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6735 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111110111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111110111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1685
#2;

verify(ir === 'b1111, "Assert 6736 : < ir !== 'b1111 >");	// Vector No: 1684
verify(op === 'b11111111, "Assert 6737 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6738 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6739 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111110111111111111111111111111111111:0:1:1011:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111110111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1686
#2;

verify(ir === 'b1011, "Assert 6740 : < ir !== 'b1011 >");	// Vector No: 1685
verify(op === 'b11111111, "Assert 6741 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6742 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6743 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111110111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111110111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1687
#2;

verify(ir === 'b1011, "Assert 6744 : < ir !== 'b1011 >");	// Vector No: 1686
verify(op === 'b11111000, "Assert 6745 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6746 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6747 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111110111111111111111111111111111111:1:1:1111:01111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111110111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1688
#2;

verify(ir === 'b1111, "Assert 6748 : < ir !== 'b1111 >");	// Vector No: 1687
verify(op === 'b01111000, "Assert 6749 : < op !== 'b01111000 >");
verify(extop === 0, "Assert 6750 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6751 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1689
#2;

verify(ir === 'b1111, "Assert 6752 : < ir !== 'b1111 >");	// Vector No: 1688
verify(op === 'b11111111, "Assert 6753 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6754 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6755 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101110011111111111111111111111111:0:1:0111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1690
#2;

verify(ir === 'b0111, "Assert 6756 : < ir !== 'b0111 >");	// Vector No: 1689
verify(op === 'b11111111, "Assert 6757 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6758 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6759 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1691
#2;

verify(ir === 'b1111, "Assert 6760 : < ir !== 'b1111 >");	// Vector No: 1690
verify(op === 'b11111000, "Assert 6761 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6762 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6763 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111101110011111111111111111111111111:1:1:1111:01110011:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111101110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1692
#2;

verify(ir === 'b1111, "Assert 6764 : < ir !== 'b1111 >");	// Vector No: 1691
verify(op === 'b01110011, "Assert 6765 : < op !== 'b01110011 >");
verify(extop === 0, "Assert 6766 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6767 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111101111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111101111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1693
#2;

verify(ir === 'b1111, "Assert 6768 : < ir !== 'b1111 >");	// Vector No: 1692
verify(op === 'b11111111, "Assert 6769 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6770 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6771 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111101111111111111111111111111111111:0:1:0111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111101111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1694
#2;

verify(ir === 'b0111, "Assert 6772 : < ir !== 'b0111 >");	// Vector No: 1693
verify(op === 'b11111111, "Assert 6773 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6774 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6775 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111101111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111101111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1695
#2;

verify(ir === 'b1011, "Assert 6776 : < ir !== 'b1011 >");	// Vector No: 1694
verify(op === 'b11111000, "Assert 6777 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6778 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6779 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111101111111111111111111111111111111:1:1:1111:01111111:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111101111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1696
#2;

verify(ir === 'b1111, "Assert 6780 : < ir !== 'b1111 >");	// Vector No: 1695
verify(op === 'b01111111, "Assert 6781 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 6782 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6783 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1697
#2;

verify(ir === 'b1111, "Assert 6784 : < ir !== 'b1111 >");	// Vector No: 1696
verify(op === 'b11111111, "Assert 6785 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6786 : < extop !== 0 >");
verify(addr === 'b11111111111111111110, "Assert 6787 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1698
#2;

verify(ir === 'b1111, "Assert 6788 : < ir !== 'b1111 >");	// Vector No: 1697
verify(op === 'b11111111, "Assert 6789 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6790 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6791 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1699
#2;

verify(ir === 'b1111, "Assert 6792 : < ir !== 'b1111 >");	// Vector No: 1698
verify(op === 'b11111000, "Assert 6793 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6794 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6795 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111111011110011111111111111111111111111:1:1:1110:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111111011110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1700
#2;

verify(ir === 'b1110, "Assert 6796 : < ir !== 'b1110 >");	// Vector No: 1699
verify(op === 'b11100000, "Assert 6797 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6798 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6799 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111011111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111110:
//------------------------

#2;
word <= 'b1111001111111111111111111111111011111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1701
#2;

verify(ir === 'b1111, "Assert 6800 : < ir !== 'b1111 >");	// Vector No: 1700
verify(op === 'b11111111, "Assert 6801 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6802 : < extop !== 1 >");
verify(addr === 'b11111111111111111110, "Assert 6803 : < addr !== 'b11111111111111111110 >");
#2;
clk <= 0;

// 1111001111111111111111111111111011111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111011111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1702
#2;

verify(ir === 'b1111, "Assert 6804 : < ir !== 'b1111 >");	// Vector No: 1701
verify(op === 'b11111111, "Assert 6805 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6806 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6807 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111011111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111011111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1703
#2;

verify(ir === 'b1011, "Assert 6808 : < ir !== 'b1011 >");	// Vector No: 1702
verify(op === 'b11111000, "Assert 6809 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6810 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6811 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111011111111111111111111111111111111:1:1:1110:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111011111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1704
#2;

verify(ir === 'b1110, "Assert 6812 : < ir !== 'b1110 >");	// Vector No: 1703
verify(op === 'b11111000, "Assert 6813 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6814 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6815 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1705
#2;

verify(ir === 'b1111, "Assert 6816 : < ir !== 'b1111 >");	// Vector No: 1704
verify(op === 'b11111111, "Assert 6817 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6818 : < extop !== 0 >");
verify(addr === 'b11111111111111111101, "Assert 6819 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1706
#2;

verify(ir === 'b1111, "Assert 6820 : < ir !== 'b1111 >");	// Vector No: 1705
verify(op === 'b11111111, "Assert 6821 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6822 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6823 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1707
#2;

verify(ir === 'b1111, "Assert 6824 : < ir !== 'b1111 >");	// Vector No: 1706
verify(op === 'b11111000, "Assert 6825 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6826 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6827 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111110111110011111111111111111111111111:1:1:1101:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111110111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1708
#2;

verify(ir === 'b1101, "Assert 6828 : < ir !== 'b1101 >");	// Vector No: 1707
verify(op === 'b11100000, "Assert 6829 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6830 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6831 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111110111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111101:
//------------------------

#2;
word <= 'b1111001111111111111111111111110111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1709
#2;

verify(ir === 'b1111, "Assert 6832 : < ir !== 'b1111 >");	// Vector No: 1708
verify(op === 'b11111111, "Assert 6833 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6834 : < extop !== 1 >");
verify(addr === 'b11111111111111111101, "Assert 6835 : < addr !== 'b11111111111111111101 >");
#2;
clk <= 0;

// 1111001111111111111111111111110111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111110111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1710
#2;

verify(ir === 'b1111, "Assert 6836 : < ir !== 'b1111 >");	// Vector No: 1709
verify(op === 'b11111111, "Assert 6837 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6838 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6839 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111110111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111110111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1711
#2;

verify(ir === 'b1011, "Assert 6840 : < ir !== 'b1011 >");	// Vector No: 1710
verify(op === 'b11111000, "Assert 6841 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6842 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6843 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111110111111111111111111111111111111111:1:1:1101:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111110111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1712
#2;

verify(ir === 'b1101, "Assert 6844 : < ir !== 'b1101 >");	// Vector No: 1711
verify(op === 'b11111000, "Assert 6845 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6846 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6847 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1713
#2;

verify(ir === 'b1111, "Assert 6848 : < ir !== 'b1111 >");	// Vector No: 1712
verify(op === 'b11111111, "Assert 6849 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6850 : < extop !== 0 >");
verify(addr === 'b11111111111111111011, "Assert 6851 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1714
#2;

verify(ir === 'b1111, "Assert 6852 : < ir !== 'b1111 >");	// Vector No: 1713
verify(op === 'b11111111, "Assert 6853 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6854 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6855 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1715
#2;

verify(ir === 'b1111, "Assert 6856 : < ir !== 'b1111 >");	// Vector No: 1714
verify(op === 'b11111000, "Assert 6857 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6858 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6859 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111101111110011111111111111111111111111:1:1:1011:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111101111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1716
#2;

verify(ir === 'b1011, "Assert 6860 : < ir !== 'b1011 >");	// Vector No: 1715
verify(op === 'b11100000, "Assert 6861 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6862 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6863 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111101111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111011:
//------------------------

#2;
word <= 'b1111001111111111111111111111101111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1717
#2;

verify(ir === 'b1111, "Assert 6864 : < ir !== 'b1111 >");	// Vector No: 1716
verify(op === 'b11111111, "Assert 6865 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6866 : < extop !== 1 >");
verify(addr === 'b11111111111111111011, "Assert 6867 : < addr !== 'b11111111111111111011 >");
#2;
clk <= 0;

// 1111001111111111111111111111101111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111101111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1718
#2;

verify(ir === 'b1111, "Assert 6868 : < ir !== 'b1111 >");	// Vector No: 1717
verify(op === 'b11111111, "Assert 6869 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6870 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6871 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111101111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111101111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1719
#2;

verify(ir === 'b1011, "Assert 6872 : < ir !== 'b1011 >");	// Vector No: 1718
verify(op === 'b11111000, "Assert 6873 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6874 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6875 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111101111111111111111111111111111111111:1:1:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111101111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1720
#2;

verify(ir === 'b1011, "Assert 6876 : < ir !== 'b1011 >");	// Vector No: 1719
verify(op === 'b11111000, "Assert 6877 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6878 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6879 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1721
#2;

verify(ir === 'b1111, "Assert 6880 : < ir !== 'b1111 >");	// Vector No: 1720
verify(op === 'b11111111, "Assert 6881 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6882 : < extop !== 0 >");
verify(addr === 'b11111111111111110111, "Assert 6883 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1722
#2;

verify(ir === 'b1111, "Assert 6884 : < ir !== 'b1111 >");	// Vector No: 1721
verify(op === 'b11111111, "Assert 6885 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6886 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6887 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1723
#2;

verify(ir === 'b1111, "Assert 6888 : < ir !== 'b1111 >");	// Vector No: 1722
verify(op === 'b11111000, "Assert 6889 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6890 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6891 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111111011111110011111111111111111111111111:1:1:0111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111111011111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1724
#2;

verify(ir === 'b0111, "Assert 6892 : < ir !== 'b0111 >");	// Vector No: 1723
verify(op === 'b11100000, "Assert 6893 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6894 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6895 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111011111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111110111:
//------------------------

#2;
word <= 'b1111001111111111111111111111011111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1725
#2;

verify(ir === 'b1111, "Assert 6896 : < ir !== 'b1111 >");	// Vector No: 1724
verify(op === 'b11111111, "Assert 6897 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6898 : < extop !== 1 >");
verify(addr === 'b11111111111111110111, "Assert 6899 : < addr !== 'b11111111111111110111 >");
#2;
clk <= 0;

// 1111001111111111111111111111011111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111011111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1726
#2;

verify(ir === 'b1111, "Assert 6900 : < ir !== 'b1111 >");	// Vector No: 1725
verify(op === 'b11111111, "Assert 6901 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6902 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6903 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111011111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111011111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1727
#2;

verify(ir === 'b1011, "Assert 6904 : < ir !== 'b1011 >");	// Vector No: 1726
verify(op === 'b11111000, "Assert 6905 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6906 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6907 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111011111111111111111111111111111111111:1:1:0111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111011111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1728
#2;

verify(ir === 'b0111, "Assert 6908 : < ir !== 'b0111 >");	// Vector No: 1727
verify(op === 'b11111000, "Assert 6909 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6910 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6911 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1729
#2;

verify(ir === 'b1111, "Assert 6912 : < ir !== 'b1111 >");	// Vector No: 1728
verify(op === 'b11111111, "Assert 6913 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6914 : < extop !== 0 >");
verify(addr === 'b11111111111111101111, "Assert 6915 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1730
#2;

verify(ir === 'b1111, "Assert 6916 : < ir !== 'b1111 >");	// Vector No: 1729
verify(op === 'b11111111, "Assert 6917 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6918 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6919 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111110:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1731
#2;

verify(ir === 'b1111, "Assert 6920 : < ir !== 'b1111 >");	// Vector No: 1730
verify(op === 'b11111000, "Assert 6921 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6922 : < extop !== 0 >");
verify(addr === 'b00000111111111111110, "Assert 6923 : < addr !== 'b00000111111111111110 >");
#2;
clk <= 0;

// 1111111111111111111111111110111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111110111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1732
#2;

verify(ir === 'b1111, "Assert 6924 : < ir !== 'b1111 >");	// Vector No: 1731
verify(op === 'b11100000, "Assert 6925 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6926 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6927 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111110111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111101111:
//------------------------

#2;
word <= 'b1111001111111111111111111110111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1733
#2;

verify(ir === 'b1111, "Assert 6928 : < ir !== 'b1111 >");	// Vector No: 1732
verify(op === 'b11111111, "Assert 6929 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6930 : < extop !== 1 >");
verify(addr === 'b11111111111111101111, "Assert 6931 : < addr !== 'b11111111111111101111 >");
#2;
clk <= 0;

// 1111001111111111111111111110111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111110111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1734
#2;

verify(ir === 'b1111, "Assert 6932 : < ir !== 'b1111 >");	// Vector No: 1733
verify(op === 'b11111111, "Assert 6933 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6934 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6935 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111110111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111110:
//------------------------

#2;
word <= 'b1111001111111111111111111110111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1735
#2;

verify(ir === 'b1011, "Assert 6936 : < ir !== 'b1011 >");	// Vector No: 1734
verify(op === 'b11111000, "Assert 6937 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6938 : < extop !== 0 >");
verify(addr === 'b00000111111111111110, "Assert 6939 : < addr !== 'b00000111111111111110 >");
#2;
clk <= 0;

// 1111001111111111111111111110111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111110111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1736
#2;

verify(ir === 'b1111, "Assert 6940 : < ir !== 'b1111 >");	// Vector No: 1735
verify(op === 'b11111000, "Assert 6941 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6942 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6943 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1737
#2;

verify(ir === 'b1111, "Assert 6944 : < ir !== 'b1111 >");	// Vector No: 1736
verify(op === 'b11111111, "Assert 6945 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6946 : < extop !== 0 >");
verify(addr === 'b11111111111111011111, "Assert 6947 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1738
#2;

verify(ir === 'b1111, "Assert 6948 : < ir !== 'b1111 >");	// Vector No: 1737
verify(op === 'b11111111, "Assert 6949 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6950 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6951 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111101:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1739
#2;

verify(ir === 'b1111, "Assert 6952 : < ir !== 'b1111 >");	// Vector No: 1738
verify(op === 'b11111000, "Assert 6953 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6954 : < extop !== 0 >");
verify(addr === 'b00000111111111111101, "Assert 6955 : < addr !== 'b00000111111111111101 >");
#2;
clk <= 0;

// 1111111111111111111111111101111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111101111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1740
#2;

verify(ir === 'b1111, "Assert 6956 : < ir !== 'b1111 >");	// Vector No: 1739
verify(op === 'b11100000, "Assert 6957 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6958 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6959 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111101111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111011111:
//------------------------

#2;
word <= 'b1111001111111111111111111101111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1741
#2;

verify(ir === 'b1111, "Assert 6960 : < ir !== 'b1111 >");	// Vector No: 1740
verify(op === 'b11111111, "Assert 6961 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6962 : < extop !== 1 >");
verify(addr === 'b11111111111111011111, "Assert 6963 : < addr !== 'b11111111111111011111 >");
#2;
clk <= 0;

// 1111001111111111111111111101111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111101111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1742
#2;

verify(ir === 'b1111, "Assert 6964 : < ir !== 'b1111 >");	// Vector No: 1741
verify(op === 'b11111111, "Assert 6965 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6966 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6967 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111101111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111101:
//------------------------

#2;
word <= 'b1111001111111111111111111101111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1743
#2;

verify(ir === 'b1011, "Assert 6968 : < ir !== 'b1011 >");	// Vector No: 1742
verify(op === 'b11111000, "Assert 6969 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6970 : < extop !== 0 >");
verify(addr === 'b00000111111111111101, "Assert 6971 : < addr !== 'b00000111111111111101 >");
#2;
clk <= 0;

// 1111001111111111111111111101111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111101111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1744
#2;

verify(ir === 'b1111, "Assert 6972 : < ir !== 'b1111 >");	// Vector No: 1743
verify(op === 'b11111000, "Assert 6973 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6974 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 6975 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1745
#2;

verify(ir === 'b1111, "Assert 6976 : < ir !== 'b1111 >");	// Vector No: 1744
verify(op === 'b11111111, "Assert 6977 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6978 : < extop !== 0 >");
verify(addr === 'b11111111111110111111, "Assert 6979 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1746
#2;

verify(ir === 'b1111, "Assert 6980 : < ir !== 'b1111 >");	// Vector No: 1745
verify(op === 'b11111111, "Assert 6981 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6982 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 6983 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111011:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1747
#2;

verify(ir === 'b1111, "Assert 6984 : < ir !== 'b1111 >");	// Vector No: 1746
verify(op === 'b11111000, "Assert 6985 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 6986 : < extop !== 0 >");
verify(addr === 'b00000111111111111011, "Assert 6987 : < addr !== 'b00000111111111111011 >");
#2;
clk <= 0;

// 1111111111111111111111111011111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111111011111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1748
#2;

verify(ir === 'b1111, "Assert 6988 : < ir !== 'b1111 >");	// Vector No: 1747
verify(op === 'b11100000, "Assert 6989 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 6990 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 6991 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111011111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111110111111:
//------------------------

#2;
word <= 'b1111001111111111111111111011111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1749
#2;

verify(ir === 'b1111, "Assert 6992 : < ir !== 'b1111 >");	// Vector No: 1748
verify(op === 'b11111111, "Assert 6993 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 6994 : < extop !== 1 >");
verify(addr === 'b11111111111110111111, "Assert 6995 : < addr !== 'b11111111111110111111 >");
#2;
clk <= 0;

// 1111001111111111111111111011111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111011111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1750
#2;

verify(ir === 'b1111, "Assert 6996 : < ir !== 'b1111 >");	// Vector No: 1749
verify(op === 'b11111111, "Assert 6997 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 6998 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 6999 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111011111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111011:
//------------------------

#2;
word <= 'b1111001111111111111111111011111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1751
#2;

verify(ir === 'b1011, "Assert 7000 : < ir !== 'b1011 >");	// Vector No: 1750
verify(op === 'b11111000, "Assert 7001 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7002 : < extop !== 0 >");
verify(addr === 'b00000111111111111011, "Assert 7003 : < addr !== 'b00000111111111111011 >");
#2;
clk <= 0;

// 1111001111111111111111111011111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111011111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1752
#2;

verify(ir === 'b1111, "Assert 7004 : < ir !== 'b1111 >");	// Vector No: 1751
verify(op === 'b11111000, "Assert 7005 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7006 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7007 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1753
#2;

verify(ir === 'b1111, "Assert 7008 : < ir !== 'b1111 >");	// Vector No: 1752
verify(op === 'b11111111, "Assert 7009 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7010 : < extop !== 0 >");
verify(addr === 'b11111111111101111111, "Assert 7011 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1754
#2;

verify(ir === 'b1111, "Assert 7012 : < ir !== 'b1111 >");	// Vector No: 1753
verify(op === 'b11111111, "Assert 7013 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7014 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7015 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111110111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1755
#2;

verify(ir === 'b1111, "Assert 7016 : < ir !== 'b1111 >");	// Vector No: 1754
verify(op === 'b11111000, "Assert 7017 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7018 : < extop !== 0 >");
verify(addr === 'b00000111111111110111, "Assert 7019 : < addr !== 'b00000111111111110111 >");
#2;
clk <= 0;

// 1111111111111111111111110111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111110111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1756
#2;

verify(ir === 'b1111, "Assert 7020 : < ir !== 'b1111 >");	// Vector No: 1755
verify(op === 'b11100000, "Assert 7021 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7022 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7023 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111110111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111101111111:
//------------------------

#2;
word <= 'b1111001111111111111111110111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1757
#2;

verify(ir === 'b1111, "Assert 7024 : < ir !== 'b1111 >");	// Vector No: 1756
verify(op === 'b11111111, "Assert 7025 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7026 : < extop !== 1 >");
verify(addr === 'b11111111111101111111, "Assert 7027 : < addr !== 'b11111111111101111111 >");
#2;
clk <= 0;

// 1111001111111111111111110111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111110111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1758
#2;

verify(ir === 'b1111, "Assert 7028 : < ir !== 'b1111 >");	// Vector No: 1757
verify(op === 'b11111111, "Assert 7029 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7030 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7031 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111110111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111110111:
//------------------------

#2;
word <= 'b1111001111111111111111110111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1759
#2;

verify(ir === 'b1011, "Assert 7032 : < ir !== 'b1011 >");	// Vector No: 1758
verify(op === 'b11111000, "Assert 7033 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7034 : < extop !== 0 >");
verify(addr === 'b00000111111111110111, "Assert 7035 : < addr !== 'b00000111111111110111 >");
#2;
clk <= 0;

// 1111001111111111111111110111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111110111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1760
#2;

verify(ir === 'b1111, "Assert 7036 : < ir !== 'b1111 >");	// Vector No: 1759
verify(op === 'b11111000, "Assert 7037 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7038 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7039 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1761
#2;

verify(ir === 'b1111, "Assert 7040 : < ir !== 'b1111 >");	// Vector No: 1760
verify(op === 'b11111111, "Assert 7041 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7042 : < extop !== 0 >");
verify(addr === 'b11111111111011111111, "Assert 7043 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1762
#2;

verify(ir === 'b1111, "Assert 7044 : < ir !== 'b1111 >");	// Vector No: 1761
verify(op === 'b11111111, "Assert 7045 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7046 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7047 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111101111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1763
#2;

verify(ir === 'b1111, "Assert 7048 : < ir !== 'b1111 >");	// Vector No: 1762
verify(op === 'b11111000, "Assert 7049 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7050 : < extop !== 0 >");
verify(addr === 'b00000111111111101111, "Assert 7051 : < addr !== 'b00000111111111101111 >");
#2;
clk <= 0;

// 1111111111111111111111101111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111101111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1764
#2;

verify(ir === 'b1111, "Assert 7052 : < ir !== 'b1111 >");	// Vector No: 1763
verify(op === 'b11100000, "Assert 7053 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7054 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7055 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111101111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111011111111:
//------------------------

#2;
word <= 'b1111001111111111111111101111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1765
#2;

verify(ir === 'b1111, "Assert 7056 : < ir !== 'b1111 >");	// Vector No: 1764
verify(op === 'b11111111, "Assert 7057 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7058 : < extop !== 1 >");
verify(addr === 'b11111111111011111111, "Assert 7059 : < addr !== 'b11111111111011111111 >");
#2;
clk <= 0;

// 1111001111111111111111101111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111101111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1766
#2;

verify(ir === 'b1111, "Assert 7060 : < ir !== 'b1111 >");	// Vector No: 1765
verify(op === 'b11111111, "Assert 7061 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7062 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7063 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111101111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111101111:
//------------------------

#2;
word <= 'b1111001111111111111111101111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1767
#2;

verify(ir === 'b1011, "Assert 7064 : < ir !== 'b1011 >");	// Vector No: 1766
verify(op === 'b11111000, "Assert 7065 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7066 : < extop !== 0 >");
verify(addr === 'b00000111111111101111, "Assert 7067 : < addr !== 'b00000111111111101111 >");
#2;
clk <= 0;

// 1111001111111111111111101111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111101111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1768
#2;

verify(ir === 'b1111, "Assert 7068 : < ir !== 'b1111 >");	// Vector No: 1767
verify(op === 'b11111000, "Assert 7069 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7070 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7071 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111110111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1769
#2;

verify(ir === 'b1111, "Assert 7072 : < ir !== 'b1111 >");	// Vector No: 1768
verify(op === 'b11111111, "Assert 7073 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7074 : < extop !== 0 >");
verify(addr === 'b11111111110111111111, "Assert 7075 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1770
#2;

verify(ir === 'b1111, "Assert 7076 : < ir !== 'b1111 >");	// Vector No: 1769
verify(op === 'b11111111, "Assert 7077 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7078 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7079 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111011111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1771
#2;

verify(ir === 'b1111, "Assert 7080 : < ir !== 'b1111 >");	// Vector No: 1770
verify(op === 'b11111000, "Assert 7081 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7082 : < extop !== 0 >");
verify(addr === 'b00000111111111011111, "Assert 7083 : < addr !== 'b00000111111111011111 >");
#2;
clk <= 0;

// 1111111111111111111111011111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111111011111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1772
#2;

verify(ir === 'b1111, "Assert 7084 : < ir !== 'b1111 >");	// Vector No: 1771
verify(op === 'b11100000, "Assert 7085 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7086 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7087 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111011111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111110111111111:
//------------------------

#2;
word <= 'b1111001111111111111111011111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1773
#2;

verify(ir === 'b1111, "Assert 7088 : < ir !== 'b1111 >");	// Vector No: 1772
verify(op === 'b11111111, "Assert 7089 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7090 : < extop !== 1 >");
verify(addr === 'b11111111110111111111, "Assert 7091 : < addr !== 'b11111111110111111111 >");
#2;
clk <= 0;

// 1111001111111111111111011111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111011111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1774
#2;

verify(ir === 'b1111, "Assert 7092 : < ir !== 'b1111 >");	// Vector No: 1773
verify(op === 'b11111111, "Assert 7093 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7094 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7095 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111011111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111011111:
//------------------------

#2;
word <= 'b1111001111111111111111011111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1775
#2;

verify(ir === 'b1011, "Assert 7096 : < ir !== 'b1011 >");	// Vector No: 1774
verify(op === 'b11111000, "Assert 7097 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7098 : < extop !== 0 >");
verify(addr === 'b00000111111111011111, "Assert 7099 : < addr !== 'b00000111111111011111 >");
#2;
clk <= 0;

// 1111001111111111111111011111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111011111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1776
#2;

verify(ir === 'b1111, "Assert 7100 : < ir !== 'b1111 >");	// Vector No: 1775
verify(op === 'b11111000, "Assert 7101 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7102 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7103 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111101111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1777
#2;

verify(ir === 'b1111, "Assert 7104 : < ir !== 'b1111 >");	// Vector No: 1776
verify(op === 'b11111111, "Assert 7105 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7106 : < extop !== 0 >");
verify(addr === 'b11111111101111111111, "Assert 7107 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1778
#2;

verify(ir === 'b1111, "Assert 7108 : < ir !== 'b1111 >");	// Vector No: 1777
verify(op === 'b11111111, "Assert 7109 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7110 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7111 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111110111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1779
#2;

verify(ir === 'b1111, "Assert 7112 : < ir !== 'b1111 >");	// Vector No: 1778
verify(op === 'b11111000, "Assert 7113 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7114 : < extop !== 0 >");
verify(addr === 'b00000111111110111111, "Assert 7115 : < addr !== 'b00000111111110111111 >");
#2;
clk <= 0;

// 1111111111111111111110111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111110111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1780
#2;

verify(ir === 'b1111, "Assert 7116 : < ir !== 'b1111 >");	// Vector No: 1779
verify(op === 'b11100000, "Assert 7117 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7118 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7119 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111110111111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111101111111111:
//------------------------

#2;
word <= 'b1111001111111111111110111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1781
#2;

verify(ir === 'b1111, "Assert 7120 : < ir !== 'b1111 >");	// Vector No: 1780
verify(op === 'b11111111, "Assert 7121 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7122 : < extop !== 1 >");
verify(addr === 'b11111111101111111111, "Assert 7123 : < addr !== 'b11111111101111111111 >");
#2;
clk <= 0;

// 1111001111111111111110111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111110111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1782
#2;

verify(ir === 'b1111, "Assert 7124 : < ir !== 'b1111 >");	// Vector No: 1781
verify(op === 'b11111111, "Assert 7125 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7126 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7127 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111110111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111110111111:
//------------------------

#2;
word <= 'b1111001111111111111110111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1783
#2;

verify(ir === 'b1011, "Assert 7128 : < ir !== 'b1011 >");	// Vector No: 1782
verify(op === 'b11111000, "Assert 7129 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7130 : < extop !== 0 >");
verify(addr === 'b00000111111110111111, "Assert 7131 : < addr !== 'b00000111111110111111 >");
#2;
clk <= 0;

// 1111001111111111111110111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111110111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1784
#2;

verify(ir === 'b1111, "Assert 7132 : < ir !== 'b1111 >");	// Vector No: 1783
verify(op === 'b11111000, "Assert 7133 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7134 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7135 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111111011111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1785
#2;

verify(ir === 'b1111, "Assert 7136 : < ir !== 'b1111 >");	// Vector No: 1784
verify(op === 'b11111111, "Assert 7137 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7138 : < extop !== 0 >");
verify(addr === 'b11111111011111111111, "Assert 7139 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1786
#2;

verify(ir === 'b1111, "Assert 7140 : < ir !== 'b1111 >");	// Vector No: 1785
verify(op === 'b11111111, "Assert 7141 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7142 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7143 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111101111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1787
#2;

verify(ir === 'b1111, "Assert 7144 : < ir !== 'b1111 >");	// Vector No: 1786
verify(op === 'b11111000, "Assert 7145 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7146 : < extop !== 0 >");
verify(addr === 'b00000111111101111111, "Assert 7147 : < addr !== 'b00000111111101111111 >");
#2;
clk <= 0;

// 1111111111111111111101111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111101111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1788
#2;

verify(ir === 'b1111, "Assert 7148 : < ir !== 'b1111 >");	// Vector No: 1787
verify(op === 'b11100000, "Assert 7149 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7150 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7151 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111101111111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111011111111111:
//------------------------

#2;
word <= 'b1111001111111111111101111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1789
#2;

verify(ir === 'b1111, "Assert 7152 : < ir !== 'b1111 >");	// Vector No: 1788
verify(op === 'b11111111, "Assert 7153 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7154 : < extop !== 1 >");
verify(addr === 'b11111111011111111111, "Assert 7155 : < addr !== 'b11111111011111111111 >");
#2;
clk <= 0;

// 1111001111111111111101111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111101111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1790
#2;

verify(ir === 'b1111, "Assert 7156 : < ir !== 'b1111 >");	// Vector No: 1789
verify(op === 'b11111111, "Assert 7157 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7158 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7159 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111101111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111101111111:
//------------------------

#2;
word <= 'b1111001111111111111101111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1791
#2;

verify(ir === 'b1011, "Assert 7160 : < ir !== 'b1011 >");	// Vector No: 1790
verify(op === 'b11111000, "Assert 7161 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7162 : < extop !== 0 >");
verify(addr === 'b00000111111101111111, "Assert 7163 : < addr !== 'b00000111111101111111 >");
#2;
clk <= 0;

// 1111001111111111111101111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111101111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1792
#2;

verify(ir === 'b1111, "Assert 7164 : < ir !== 'b1111 >");	// Vector No: 1791
verify(op === 'b11111000, "Assert 7165 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7166 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7167 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111110111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1793
#2;

verify(ir === 'b1111, "Assert 7168 : < ir !== 'b1111 >");	// Vector No: 1792
verify(op === 'b11111111, "Assert 7169 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7170 : < extop !== 0 >");
verify(addr === 'b11111110111111111111, "Assert 7171 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1794
#2;

verify(ir === 'b1111, "Assert 7172 : < ir !== 'b1111 >");	// Vector No: 1793
verify(op === 'b11111111, "Assert 7173 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7174 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7175 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111011111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1795
#2;

verify(ir === 'b1111, "Assert 7176 : < ir !== 'b1111 >");	// Vector No: 1794
verify(op === 'b11111000, "Assert 7177 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7178 : < extop !== 0 >");
verify(addr === 'b00000111111011111111, "Assert 7179 : < addr !== 'b00000111111011111111 >");
#2;
clk <= 0;

// 1111111111111111111011111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111111011111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1796
#2;

verify(ir === 'b1111, "Assert 7180 : < ir !== 'b1111 >");	// Vector No: 1795
verify(op === 'b11100000, "Assert 7181 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7182 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7183 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111011111111111111111111111111111111111111111111:0:0:1111:11111110:1:11111110111111111111:
//------------------------

#2;
word <= 'b1111001111111111111011111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1797
#2;

verify(ir === 'b1111, "Assert 7184 : < ir !== 'b1111 >");	// Vector No: 1796
verify(op === 'b11111110, "Assert 7185 : < op !== 'b11111110 >");
verify(extop === 1, "Assert 7186 : < extop !== 1 >");
verify(addr === 'b11111110111111111111, "Assert 7187 : < addr !== 'b11111110111111111111 >");
#2;
clk <= 0;

// 1111001111111111111011111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111011111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1798
#2;

verify(ir === 'b1111, "Assert 7188 : < ir !== 'b1111 >");	// Vector No: 1797
verify(op === 'b11111111, "Assert 7189 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7190 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7191 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111011111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111011111111:
//------------------------

#2;
word <= 'b1111001111111111111011111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1799
#2;

verify(ir === 'b1011, "Assert 7192 : < ir !== 'b1011 >");	// Vector No: 1798
verify(op === 'b11111000, "Assert 7193 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7194 : < extop !== 0 >");
verify(addr === 'b00000111111011111111, "Assert 7195 : < addr !== 'b00000111111011111111 >");
#2;
clk <= 0;

// 1111001111111111111011111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111011111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1800
#2;

verify(ir === 'b1111, "Assert 7196 : < ir !== 'b1111 >");	// Vector No: 1799
verify(op === 'b11111000, "Assert 7197 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7198 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7199 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111101111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1801
#2;

verify(ir === 'b1111, "Assert 7200 : < ir !== 'b1111 >");	// Vector No: 1800
verify(op === 'b11111111, "Assert 7201 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7202 : < extop !== 0 >");
verify(addr === 'b11111101111111111111, "Assert 7203 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1802
#2;

verify(ir === 'b1111, "Assert 7204 : < ir !== 'b1111 >");	// Vector No: 1801
verify(op === 'b11111111, "Assert 7205 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7206 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7207 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111110111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1803
#2;

verify(ir === 'b1111, "Assert 7208 : < ir !== 'b1111 >");	// Vector No: 1802
verify(op === 'b11111000, "Assert 7209 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7210 : < extop !== 0 >");
verify(addr === 'b00000111110111111111, "Assert 7211 : < addr !== 'b00000111110111111111 >");
#2;
clk <= 0;

// 1111111111111111110111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111110111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1804
#2;

verify(ir === 'b1111, "Assert 7212 : < ir !== 'b1111 >");	// Vector No: 1803
verify(op === 'b11100000, "Assert 7213 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7214 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7215 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111110111111111111111111111111111111111111111111111:0:0:1111:11111101:1:11111101111111111111:
//------------------------

#2;
word <= 'b1111001111111111110111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1805
#2;

verify(ir === 'b1111, "Assert 7216 : < ir !== 'b1111 >");	// Vector No: 1804
verify(op === 'b11111101, "Assert 7217 : < op !== 'b11111101 >");
verify(extop === 1, "Assert 7218 : < extop !== 1 >");
verify(addr === 'b11111101111111111111, "Assert 7219 : < addr !== 'b11111101111111111111 >");
#2;
clk <= 0;

// 1111001111111111110111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111110111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1806
#2;

verify(ir === 'b1111, "Assert 7220 : < ir !== 'b1111 >");	// Vector No: 1805
verify(op === 'b11111111, "Assert 7221 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7222 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7223 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111110111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111110111111111:
//------------------------

#2;
word <= 'b1111001111111111110111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1807
#2;

verify(ir === 'b1011, "Assert 7224 : < ir !== 'b1011 >");	// Vector No: 1806
verify(op === 'b11111000, "Assert 7225 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7226 : < extop !== 0 >");
verify(addr === 'b00000111110111111111, "Assert 7227 : < addr !== 'b00000111110111111111 >");
#2;
clk <= 0;

// 1111001111111111110111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111110111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1808
#2;

verify(ir === 'b1111, "Assert 7228 : < ir !== 'b1111 >");	// Vector No: 1807
verify(op === 'b11111000, "Assert 7229 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7230 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7231 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11111011111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1809
#2;

verify(ir === 'b1111, "Assert 7232 : < ir !== 'b1111 >");	// Vector No: 1808
verify(op === 'b11111111, "Assert 7233 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7234 : < extop !== 0 >");
verify(addr === 'b11111011111111111111, "Assert 7235 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1810
#2;

verify(ir === 'b1111, "Assert 7236 : < ir !== 'b1111 >");	// Vector No: 1809
verify(op === 'b11111111, "Assert 7237 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7238 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7239 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111101111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1811
#2;

verify(ir === 'b1111, "Assert 7240 : < ir !== 'b1111 >");	// Vector No: 1810
verify(op === 'b11111000, "Assert 7241 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7242 : < extop !== 0 >");
verify(addr === 'b00000111101111111111, "Assert 7243 : < addr !== 'b00000111101111111111 >");
#2;
clk <= 0;

// 1111111111111111101111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111101111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1812
#2;

verify(ir === 'b1111, "Assert 7244 : < ir !== 'b1111 >");	// Vector No: 1811
verify(op === 'b11100000, "Assert 7245 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7246 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7247 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111101111111111111111111111111111111111111111111111:0:0:1111:11111011:1:11111011111111111111:
//------------------------

#2;
word <= 'b1111001111111111101111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1813
#2;

verify(ir === 'b1111, "Assert 7248 : < ir !== 'b1111 >");	// Vector No: 1812
verify(op === 'b11111011, "Assert 7249 : < op !== 'b11111011 >");
verify(extop === 1, "Assert 7250 : < extop !== 1 >");
verify(addr === 'b11111011111111111111, "Assert 7251 : < addr !== 'b11111011111111111111 >");
#2;
clk <= 0;

// 1111001111111111101111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111101111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1814
#2;

verify(ir === 'b1111, "Assert 7252 : < ir !== 'b1111 >");	// Vector No: 1813
verify(op === 'b11111111, "Assert 7253 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7254 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7255 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111101111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111101111111111:
//------------------------

#2;
word <= 'b1111001111111111101111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1815
#2;

verify(ir === 'b1011, "Assert 7256 : < ir !== 'b1011 >");	// Vector No: 1814
verify(op === 'b11111000, "Assert 7257 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7258 : < extop !== 0 >");
verify(addr === 'b00000111101111111111, "Assert 7259 : < addr !== 'b00000111101111111111 >");
#2;
clk <= 0;

// 1111001111111111101111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111101111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1816
#2;

verify(ir === 'b1111, "Assert 7260 : < ir !== 'b1111 >");	// Vector No: 1815
verify(op === 'b11111000, "Assert 7261 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7262 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7263 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11110111111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1817
#2;

verify(ir === 'b1111, "Assert 7264 : < ir !== 'b1111 >");	// Vector No: 1816
verify(op === 'b11111111, "Assert 7265 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7266 : < extop !== 0 >");
verify(addr === 'b11110111111111111111, "Assert 7267 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1818
#2;

verify(ir === 'b1111, "Assert 7268 : < ir !== 'b1111 >");	// Vector No: 1817
verify(op === 'b11111111, "Assert 7269 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7270 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7271 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111011111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1819
#2;

verify(ir === 'b1111, "Assert 7272 : < ir !== 'b1111 >");	// Vector No: 1818
verify(op === 'b11111000, "Assert 7273 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7274 : < extop !== 0 >");
verify(addr === 'b00000111011111111111, "Assert 7275 : < addr !== 'b00000111011111111111 >");
#2;
clk <= 0;

// 1111111111111111011111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111111011111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1820
#2;

verify(ir === 'b1111, "Assert 7276 : < ir !== 'b1111 >");	// Vector No: 1819
verify(op === 'b11100000, "Assert 7277 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7278 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7279 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111011111111111111111111111111111111111111111111111:0:0:1111:11110111:1:11110111111111111111:
//------------------------

#2;
word <= 'b1111001111111111011111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1821
#2;

verify(ir === 'b1111, "Assert 7280 : < ir !== 'b1111 >");	// Vector No: 1820
verify(op === 'b11110111, "Assert 7281 : < op !== 'b11110111 >");
verify(extop === 1, "Assert 7282 : < extop !== 1 >");
verify(addr === 'b11110111111111111111, "Assert 7283 : < addr !== 'b11110111111111111111 >");
#2;
clk <= 0;

// 1111001111111111011111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111011111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1822
#2;

verify(ir === 'b1111, "Assert 7284 : < ir !== 'b1111 >");	// Vector No: 1821
verify(op === 'b11111111, "Assert 7285 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7286 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7287 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111011111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111011111111111:
//------------------------

#2;
word <= 'b1111001111111111011111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1823
#2;

verify(ir === 'b1011, "Assert 7288 : < ir !== 'b1011 >");	// Vector No: 1822
verify(op === 'b11111000, "Assert 7289 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7290 : < extop !== 0 >");
verify(addr === 'b00000111011111111111, "Assert 7291 : < addr !== 'b00000111011111111111 >");
#2;
clk <= 0;

// 1111001111111111011111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111011111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1824
#2;

verify(ir === 'b1111, "Assert 7292 : < ir !== 'b1111 >");	// Vector No: 1823
verify(op === 'b11111000, "Assert 7293 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7294 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7295 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11101111111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1825
#2;

verify(ir === 'b1111, "Assert 7296 : < ir !== 'b1111 >");	// Vector No: 1824
verify(op === 'b11111111, "Assert 7297 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7298 : < extop !== 0 >");
verify(addr === 'b11101111111111111111, "Assert 7299 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1826
#2;

verify(ir === 'b1111, "Assert 7300 : < ir !== 'b1111 >");	// Vector No: 1825
verify(op === 'b11111111, "Assert 7301 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7302 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7303 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000110111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1827
#2;

verify(ir === 'b1111, "Assert 7304 : < ir !== 'b1111 >");	// Vector No: 1826
verify(op === 'b11111000, "Assert 7305 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7306 : < extop !== 0 >");
verify(addr === 'b00000110111111111111, "Assert 7307 : < addr !== 'b00000110111111111111 >");
#2;
clk <= 0;

// 1111111111111110111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111110111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1828
#2;

verify(ir === 'b1111, "Assert 7308 : < ir !== 'b1111 >");	// Vector No: 1827
verify(op === 'b11100000, "Assert 7309 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7310 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7311 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111110111111111111111111111111111111111111111111111111:0:0:1111:11101111:1:11101111111111111111:
//------------------------

#2;
word <= 'b1111001111111110111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1829
#2;

verify(ir === 'b1111, "Assert 7312 : < ir !== 'b1111 >");	// Vector No: 1828
verify(op === 'b11101111, "Assert 7313 : < op !== 'b11101111 >");
verify(extop === 1, "Assert 7314 : < extop !== 1 >");
verify(addr === 'b11101111111111111111, "Assert 7315 : < addr !== 'b11101111111111111111 >");
#2;
clk <= 0;

// 1111001111111110111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111110111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1830
#2;

verify(ir === 'b1111, "Assert 7316 : < ir !== 'b1111 >");	// Vector No: 1829
verify(op === 'b11111111, "Assert 7317 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7318 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7319 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111110111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000110111111111111:
//------------------------

#2;
word <= 'b1111001111111110111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1831
#2;

verify(ir === 'b1011, "Assert 7320 : < ir !== 'b1011 >");	// Vector No: 1830
verify(op === 'b11111000, "Assert 7321 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7322 : < extop !== 0 >");
verify(addr === 'b00000110111111111111, "Assert 7323 : < addr !== 'b00000110111111111111 >");
#2;
clk <= 0;

// 1111001111111110111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111110111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1832
#2;

verify(ir === 'b1111, "Assert 7324 : < ir !== 'b1111 >");	// Vector No: 1831
verify(op === 'b11111000, "Assert 7325 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7326 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7327 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111110011111111111111111111111111:0:0:1111:11111111:0:11011111111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1833
#2;

verify(ir === 'b1111, "Assert 7328 : < ir !== 'b1111 >");	// Vector No: 1832
verify(op === 'b11111111, "Assert 7329 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7330 : < extop !== 0 >");
verify(addr === 'b11011111111111111111, "Assert 7331 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1834
#2;

verify(ir === 'b1111, "Assert 7332 : < ir !== 'b1111 >");	// Vector No: 1833
verify(op === 'b11111111, "Assert 7333 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7334 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7335 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000101111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1835
#2;

verify(ir === 'b1111, "Assert 7336 : < ir !== 'b1111 >");	// Vector No: 1834
verify(op === 'b11111000, "Assert 7337 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7338 : < extop !== 0 >");
verify(addr === 'b00000101111111111111, "Assert 7339 : < addr !== 'b00000101111111111111 >");
#2;
clk <= 0;

// 1111111111111101111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111101111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1836
#2;

verify(ir === 'b1111, "Assert 7340 : < ir !== 'b1111 >");	// Vector No: 1835
verify(op === 'b11100000, "Assert 7341 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7342 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7343 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111101111111111111111111111111111111111111111111111111:0:0:1111:11011111:1:11011111111111111111:
//------------------------

#2;
word <= 'b1111001111111101111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1837
#2;

verify(ir === 'b1111, "Assert 7344 : < ir !== 'b1111 >");	// Vector No: 1836
verify(op === 'b11011111, "Assert 7345 : < op !== 'b11011111 >");
verify(extop === 1, "Assert 7346 : < extop !== 1 >");
verify(addr === 'b11011111111111111111, "Assert 7347 : < addr !== 'b11011111111111111111 >");
#2;
clk <= 0;

// 1111001111111101111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111101111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1838
#2;

verify(ir === 'b1111, "Assert 7348 : < ir !== 'b1111 >");	// Vector No: 1837
verify(op === 'b11111111, "Assert 7349 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7350 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7351 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111101111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000101111111111111:
//------------------------

#2;
word <= 'b1111001111111101111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1839
#2;

verify(ir === 'b1011, "Assert 7352 : < ir !== 'b1011 >");	// Vector No: 1838
verify(op === 'b11111000, "Assert 7353 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7354 : < extop !== 0 >");
verify(addr === 'b00000101111111111111, "Assert 7355 : < addr !== 'b00000101111111111111 >");
#2;
clk <= 0;

// 1111001111111101111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111101111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1840
#2;

verify(ir === 'b1111, "Assert 7356 : < ir !== 'b1111 >");	// Vector No: 1839
verify(op === 'b11111000, "Assert 7357 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7358 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7359 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111110011111111111111111111111111:0:0:1111:11111111:0:10111111111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1841
#2;

verify(ir === 'b1111, "Assert 7360 : < ir !== 'b1111 >");	// Vector No: 1840
verify(op === 'b11111111, "Assert 7361 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7362 : < extop !== 0 >");
verify(addr === 'b10111111111111111111, "Assert 7363 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1842
#2;

verify(ir === 'b1111, "Assert 7364 : < ir !== 'b1111 >");	// Vector No: 1841
verify(op === 'b11111111, "Assert 7365 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7366 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7367 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1843
#2;

verify(ir === 'b1111, "Assert 7368 : < ir !== 'b1111 >");	// Vector No: 1842
verify(op === 'b11111000, "Assert 7369 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7370 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7371 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111111111011111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111111011111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1844
#2;

verify(ir === 'b1111, "Assert 7372 : < ir !== 'b1111 >");	// Vector No: 1843
verify(op === 'b11100000, "Assert 7373 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7374 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7375 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111011111111111111111111111111111111111111111111111111:0:0:1111:10111111:1:10111111111111111111:
//------------------------

#2;
word <= 'b1111001111111011111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1845
#2;

verify(ir === 'b1111, "Assert 7376 : < ir !== 'b1111 >");	// Vector No: 1844
verify(op === 'b10111111, "Assert 7377 : < op !== 'b10111111 >");
verify(extop === 1, "Assert 7378 : < extop !== 1 >");
verify(addr === 'b10111111111111111111, "Assert 7379 : < addr !== 'b10111111111111111111 >");
#2;
clk <= 0;

// 1111001111111011111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111011111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1846
#2;

verify(ir === 'b1111, "Assert 7380 : < ir !== 'b1111 >");	// Vector No: 1845
verify(op === 'b11111111, "Assert 7381 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7382 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7383 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111011111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111001111111011111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1847
#2;

verify(ir === 'b1011, "Assert 7384 : < ir !== 'b1011 >");	// Vector No: 1846
verify(op === 'b11111000, "Assert 7385 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7386 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7387 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111011111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111011111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1848
#2;

verify(ir === 'b1111, "Assert 7388 : < ir !== 'b1111 >");	// Vector No: 1847
verify(op === 'b11111000, "Assert 7389 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7390 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7391 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111110011111111111111111111111111:0:0:1111:11111111:0:01111111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1849
#2;

verify(ir === 'b1111, "Assert 7392 : < ir !== 'b1111 >");	// Vector No: 1848
verify(op === 'b11111111, "Assert 7393 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7394 : < extop !== 0 >");
verify(addr === 'b01111111111111111111, "Assert 7395 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1850
#2;

verify(ir === 'b1111, "Assert 7396 : < ir !== 'b1111 >");	// Vector No: 1849
verify(op === 'b11111111, "Assert 7397 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7398 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7399 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111110011111111111111111111111111:1:0:1111:11110000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1851
#2;

verify(ir === 'b1111, "Assert 7400 : < ir !== 'b1111 >");	// Vector No: 1850
verify(op === 'b11110000, "Assert 7401 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 7402 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7403 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111110111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111110111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1852
#2;

verify(ir === 'b1111, "Assert 7404 : < ir !== 'b1111 >");	// Vector No: 1851
verify(op === 'b11100000, "Assert 7405 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7406 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7407 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111110111111111111111111111111111111111111111111111111111:0:0:1111:01111111:1:01111111111111111111:
//------------------------

#2;
word <= 'b1111001111110111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1853
#2;

verify(ir === 'b1111, "Assert 7408 : < ir !== 'b1111 >");	// Vector No: 1852
verify(op === 'b01111111, "Assert 7409 : < op !== 'b01111111 >");
verify(extop === 1, "Assert 7410 : < extop !== 1 >");
verify(addr === 'b01111111111111111111, "Assert 7411 : < addr !== 'b01111111111111111111 >");
#2;
clk <= 0;

// 1111001111110111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111110111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1854
#2;

verify(ir === 'b1111, "Assert 7412 : < ir !== 'b1111 >");	// Vector No: 1853
verify(op === 'b11111111, "Assert 7413 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7414 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7415 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111110111111111111111111111111111111111111111111111111111:1:0:1011:11110000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111110111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1855
#2;

verify(ir === 'b1011, "Assert 7416 : < ir !== 'b1011 >");	// Vector No: 1854
verify(op === 'b11110000, "Assert 7417 : < op !== 'b11110000 >");
verify(extop === 0, "Assert 7418 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7419 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111110111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111110111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1856
#2;

verify(ir === 'b1111, "Assert 7420 : < ir !== 'b1111 >");	// Vector No: 1855
verify(op === 'b11111000, "Assert 7421 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7422 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7423 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111110011111111111111111111111111:0:0:1111:11111110:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1857
#2;

verify(ir === 'b1111, "Assert 7424 : < ir !== 'b1111 >");	// Vector No: 1856
verify(op === 'b11111110, "Assert 7425 : < op !== 'b11111110 >");
verify(extop === 0, "Assert 7426 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7427 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1858
#2;

verify(ir === 'b1111, "Assert 7428 : < ir !== 'b1111 >");	// Vector No: 1857
verify(op === 'b11111111, "Assert 7429 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7430 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7431 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111110011111111111111111111111111:1:0:1111:11101000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1859
#2;

verify(ir === 'b1111, "Assert 7432 : < ir !== 'b1111 >");	// Vector No: 1858
verify(op === 'b11101000, "Assert 7433 : < op !== 'b11101000 >");
verify(extop === 0, "Assert 7434 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7435 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111101111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111101111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1860
#2;

verify(ir === 'b1111, "Assert 7436 : < ir !== 'b1111 >");	// Vector No: 1859
verify(op === 'b11100000, "Assert 7437 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7438 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7439 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111111:0:0:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1861
#2;

verify(ir === 'b1111, "Assert 7440 : < ir !== 'b1111 >");	// Vector No: 1860
verify(op === 'b11111111, "Assert 7441 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7442 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7443 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1862
#2;

verify(ir === 'b1111, "Assert 7444 : < ir !== 'b1111 >");	// Vector No: 1861
verify(op === 'b11111111, "Assert 7445 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7446 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7447 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1863
#2;

verify(ir === 'b1011, "Assert 7448 : < ir !== 'b1011 >");	// Vector No: 1862
verify(op === 'b11111000, "Assert 7449 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7450 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7451 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111001111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1864
#2;

verify(ir === 'b1111, "Assert 7452 : < ir !== 'b1111 >");	// Vector No: 1863
verify(op === 'b11111000, "Assert 7453 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7454 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7455 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111110011111111111111111111111111:0:0:1111:11111101:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1865
#2;

verify(ir === 'b1111, "Assert 7456 : < ir !== 'b1111 >");	// Vector No: 1864
verify(op === 'b11111101, "Assert 7457 : < op !== 'b11111101 >");
verify(extop === 0, "Assert 7458 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7459 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1866
#2;

verify(ir === 'b1111, "Assert 7460 : < ir !== 'b1111 >");	// Vector No: 1865
verify(op === 'b11111111, "Assert 7461 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7462 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7463 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111110011111111111111111111111111:1:0:1111:11011000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1867
#2;

verify(ir === 'b1111, "Assert 7464 : < ir !== 'b1111 >");	// Vector No: 1866
verify(op === 'b11011000, "Assert 7465 : < op !== 'b11011000 >");
verify(extop === 0, "Assert 7466 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7467 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111111011111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111111011111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1868
#2;

verify(ir === 'b1111, "Assert 7468 : < ir !== 'b1111 >");	// Vector No: 1867
verify(op === 'b11100000, "Assert 7469 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7470 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7471 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111110011111111111111111111111111:0:0:1111:11111011:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1869
#2;

verify(ir === 'b1111, "Assert 7472 : < ir !== 'b1111 >");	// Vector No: 1868
verify(op === 'b11111011, "Assert 7473 : < op !== 'b11111011 >");
verify(extop === 0, "Assert 7474 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7475 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1870
#2;

verify(ir === 'b1111, "Assert 7476 : < ir !== 'b1111 >");	// Vector No: 1869
verify(op === 'b11111111, "Assert 7477 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7478 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7479 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111110011111111111111111111111111:1:0:1111:10111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1871
#2;

verify(ir === 'b1111, "Assert 7480 : < ir !== 'b1111 >");	// Vector No: 1870
verify(op === 'b10111000, "Assert 7481 : < op !== 'b10111000 >");
verify(extop === 0, "Assert 7482 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7483 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111110111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111110111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1872
#2;

verify(ir === 'b1111, "Assert 7484 : < ir !== 'b1111 >");	// Vector No: 1871
verify(op === 'b11100000, "Assert 7485 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7486 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7487 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111110011111111111111111111111111:0:0:1111:11110111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1873
#2;

verify(ir === 'b1111, "Assert 7488 : < ir !== 'b1111 >");	// Vector No: 1872
verify(op === 'b11110111, "Assert 7489 : < op !== 'b11110111 >");
verify(extop === 0, "Assert 7490 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7491 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1874
#2;

verify(ir === 'b1111, "Assert 7492 : < ir !== 'b1111 >");	// Vector No: 1873
verify(op === 'b11111111, "Assert 7493 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7494 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7495 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111110011111111111111111111111111:1:0:1111:01111111:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1875
#2;

verify(ir === 'b1111, "Assert 7496 : < ir !== 'b1111 >");	// Vector No: 1874
verify(op === 'b01111111, "Assert 7497 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 7498 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7499 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111101111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111101111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1876
#2;

verify(ir === 'b1111, "Assert 7500 : < ir !== 'b1111 >");	// Vector No: 1875
verify(op === 'b11100000, "Assert 7501 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7502 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7503 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111110011111111111111111111111111:0:0:1111:11101111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1877
#2;

verify(ir === 'b1111, "Assert 7504 : < ir !== 'b1111 >");	// Vector No: 1876
verify(op === 'b11101111, "Assert 7505 : < op !== 'b11101111 >");
verify(extop === 0, "Assert 7506 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7507 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1878
#2;

verify(ir === 'b1111, "Assert 7508 : < ir !== 'b1111 >");	// Vector No: 1877
verify(op === 'b11111111, "Assert 7509 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7510 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7511 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111110011111111111111111111111111:1:0:1110:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1879
#2;

verify(ir === 'b1110, "Assert 7512 : < ir !== 'b1110 >");	// Vector No: 1878
verify(op === 'b11111000, "Assert 7513 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7514 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7515 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111111011111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111111011111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1880
#2;

verify(ir === 'b1111, "Assert 7516 : < ir !== 'b1111 >");	// Vector No: 1879
verify(op === 'b11100000, "Assert 7517 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7518 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7519 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111110011111111111111111111111111:0:0:1111:11011111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1881
#2;

verify(ir === 'b1111, "Assert 7520 : < ir !== 'b1111 >");	// Vector No: 1880
verify(op === 'b11011111, "Assert 7521 : < op !== 'b11011111 >");
verify(extop === 0, "Assert 7522 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7523 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1882
#2;

verify(ir === 'b1111, "Assert 7524 : < ir !== 'b1111 >");	// Vector No: 1881
verify(op === 'b11111111, "Assert 7525 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7526 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7527 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111110011111111111111111111111111:1:0:1101:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1883
#2;

verify(ir === 'b1101, "Assert 7528 : < ir !== 'b1101 >");	// Vector No: 1882
verify(op === 'b11111000, "Assert 7529 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7530 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7531 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111110111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111110111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1884
#2;

verify(ir === 'b1111, "Assert 7532 : < ir !== 'b1111 >");	// Vector No: 1883
verify(op === 'b11100000, "Assert 7533 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7534 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7535 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111110011111111111111111111111111:0:0:1111:10111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1885
#2;

verify(ir === 'b1111, "Assert 7536 : < ir !== 'b1111 >");	// Vector No: 1884
verify(op === 'b10111111, "Assert 7537 : < op !== 'b10111111 >");
verify(extop === 0, "Assert 7538 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7539 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1886
#2;

verify(ir === 'b1111, "Assert 7540 : < ir !== 'b1111 >");	// Vector No: 1885
verify(op === 'b11111111, "Assert 7541 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7542 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7543 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111110011111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1887
#2;

verify(ir === 'b1011, "Assert 7544 : < ir !== 'b1011 >");	// Vector No: 1886
verify(op === 'b11111000, "Assert 7545 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7546 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7547 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111101111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111101111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1888
#2;

verify(ir === 'b1111, "Assert 7548 : < ir !== 'b1111 >");	// Vector No: 1887
verify(op === 'b11100000, "Assert 7549 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7550 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7551 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111110011111111111111111111111111:0:0:1111:01111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1889
#2;

verify(ir === 'b1111, "Assert 7552 : < ir !== 'b1111 >");	// Vector No: 1888
verify(op === 'b01111111, "Assert 7553 : < op !== 'b01111111 >");
verify(extop === 0, "Assert 7554 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7555 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1890
#2;

verify(ir === 'b1111, "Assert 7556 : < ir !== 'b1111 >");	// Vector No: 1889
verify(op === 'b11111111, "Assert 7557 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7558 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7559 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1891
#2;

verify(ir === 'b1111, "Assert 7560 : < ir !== 'b1111 >");	// Vector No: 1890
verify(op === 'b11111000, "Assert 7561 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7562 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7563 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1111011111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1111011111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1892
#2;

verify(ir === 'b1111, "Assert 7564 : < ir !== 'b1111 >");	// Vector No: 1891
verify(op === 'b11100000, "Assert 7565 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7566 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7567 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111110011111111111111111111111111:0:0:1110:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1893
#2;

verify(ir === 'b1110, "Assert 7568 : < ir !== 'b1110 >");	// Vector No: 1892
verify(op === 'b11111111, "Assert 7569 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7570 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7571 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1894
#2;

verify(ir === 'b1111, "Assert 7572 : < ir !== 'b1111 >");	// Vector No: 1893
verify(op === 'b11111111, "Assert 7573 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7574 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7575 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1895
#2;

verify(ir === 'b1111, "Assert 7576 : < ir !== 'b1111 >");	// Vector No: 1894
verify(op === 'b11111000, "Assert 7577 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7578 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7579 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1110111111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1110111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1896
#2;

verify(ir === 'b1111, "Assert 7580 : < ir !== 'b1111 >");	// Vector No: 1895
verify(op === 'b11100000, "Assert 7581 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7582 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7583 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1110001111111111111111111111111111111111111111111111111111111111:0:0:1110:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1110001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1897
#2;

verify(ir === 'b1110, "Assert 7584 : < ir !== 'b1110 >");	// Vector No: 1896
verify(op === 'b11111111, "Assert 7585 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7586 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7587 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110001111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1110001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1898
#2;

verify(ir === 'b1111, "Assert 7588 : < ir !== 'b1111 >");	// Vector No: 1897
verify(op === 'b11111111, "Assert 7589 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7590 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7591 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1110001111111111111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1110001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1899
#2;

verify(ir === 'b1011, "Assert 7592 : < ir !== 'b1011 >");	// Vector No: 1898
verify(op === 'b11111000, "Assert 7593 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7594 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7595 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1110001111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1110001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1900
#2;

verify(ir === 'b1111, "Assert 7596 : < ir !== 'b1111 >");	// Vector No: 1899
verify(op === 'b11111000, "Assert 7597 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7598 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7599 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111110011111111111111111111111111:0:0:1101:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1901
#2;

verify(ir === 'b1101, "Assert 7600 : < ir !== 'b1101 >");	// Vector No: 1900
verify(op === 'b11111111, "Assert 7601 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7602 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7603 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1902
#2;

verify(ir === 'b1111, "Assert 7604 : < ir !== 'b1111 >");	// Vector No: 1901
verify(op === 'b11111111, "Assert 7605 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7606 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7607 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1903
#2;

verify(ir === 'b1111, "Assert 7608 : < ir !== 'b1111 >");	// Vector No: 1902
verify(op === 'b11111000, "Assert 7609 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7610 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7611 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1101111111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1101111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1904
#2;

verify(ir === 'b1111, "Assert 7612 : < ir !== 'b1111 >");	// Vector No: 1903
verify(op === 'b11100000, "Assert 7613 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7614 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7615 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1101001111111111111111111111111111111111111111111111111111111111:0:0:1101:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1101001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1905
#2;

verify(ir === 'b1101, "Assert 7616 : < ir !== 'b1101 >");	// Vector No: 1904
verify(op === 'b11111111, "Assert 7617 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7618 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7619 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101001111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1101001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1906
#2;

verify(ir === 'b1111, "Assert 7620 : < ir !== 'b1111 >");	// Vector No: 1905
verify(op === 'b11111111, "Assert 7621 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7622 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7623 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1101001111111111111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1101001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1907
#2;

verify(ir === 'b1011, "Assert 7624 : < ir !== 'b1011 >");	// Vector No: 1906
verify(op === 'b11111000, "Assert 7625 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7626 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7627 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1101001111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1101001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1908
#2;

verify(ir === 'b1111, "Assert 7628 : < ir !== 'b1111 >");	// Vector No: 1907
verify(op === 'b11111000, "Assert 7629 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7630 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7631 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111110011111111111111111111111111:0:0:1011:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1909
#2;

verify(ir === 'b1011, "Assert 7632 : < ir !== 'b1011 >");	// Vector No: 1908
verify(op === 'b11111111, "Assert 7633 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7634 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7635 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1910
#2;

verify(ir === 'b1111, "Assert 7636 : < ir !== 'b1111 >");	// Vector No: 1909
verify(op === 'b11111111, "Assert 7637 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7638 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7639 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111110011111111111111111111111111:1:0:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1911
#2;

verify(ir === 'b1111, "Assert 7640 : < ir !== 'b1111 >");	// Vector No: 1910
verify(op === 'b11111000, "Assert 7641 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7642 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7643 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1011111111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b1011111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1912
#2;

verify(ir === 'b1111, "Assert 7644 : < ir !== 'b1111 >");	// Vector No: 1911
verify(op === 'b11100000, "Assert 7645 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7646 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7647 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 1011001111111111111111111111111111111111111111111111111111111111:0:0:1011:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b1011001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1913
#2;

verify(ir === 'b1011, "Assert 7648 : < ir !== 'b1011 >");	// Vector No: 1912
verify(op === 'b11111111, "Assert 7649 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7650 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7651 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011001111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b1011001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1914
#2;

verify(ir === 'b1111, "Assert 7652 : < ir !== 'b1111 >");	// Vector No: 1913
verify(op === 'b11111111, "Assert 7653 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7654 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7655 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 1011001111111111111111111111111111111111111111111111111111111111:1:0:1011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1011001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1915
#2;

verify(ir === 'b1011, "Assert 7656 : < ir !== 'b1011 >");	// Vector No: 1914
verify(op === 'b11111000, "Assert 7657 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7658 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7659 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 1011001111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b1011001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1916
#2;

verify(ir === 'b1111, "Assert 7660 : < ir !== 'b1111 >");	// Vector No: 1915
verify(op === 'b11111000, "Assert 7661 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7662 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7663 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111110011111111111111111111111111:0:0:0111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1917
#2;

verify(ir === 'b0111, "Assert 7664 : < ir !== 'b0111 >");	// Vector No: 1916
verify(op === 'b11111111, "Assert 7665 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7666 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7667 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111110011111111111111111111111111:0:1:1111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111110011111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1918
#2;

verify(ir === 'b1111, "Assert 7668 : < ir !== 'b1111 >");	// Vector No: 1917
verify(op === 'b11111111, "Assert 7669 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7670 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7671 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111110011111111111111111111111111:1:0:0111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1919
#2;

verify(ir === 'b0111, "Assert 7672 : < ir !== 'b0111 >");	// Vector No: 1918
verify(op === 'b11111000, "Assert 7673 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7674 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7675 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0111111111111111111111111111111111110011111111111111111111111111:1:1:1111:11100000:0:00000011111111111111:
//------------------------

#2;
word <= 'b0111111111111111111111111111111111110011111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1920
#2;

verify(ir === 'b1111, "Assert 7676 : < ir !== 'b1111 >");	// Vector No: 1919
verify(op === 'b11100000, "Assert 7677 : < op !== 'b11100000 >");
verify(extop === 0, "Assert 7678 : < extop !== 0 >");
verify(addr === 'b00000011111111111111, "Assert 7679 : < addr !== 'b00000011111111111111 >");
#2;
clk <= 0;

// 0111001111111111111111111111111111111111111111111111111111111111:0:0:0111:11111111:1:11111111111111111111:
//------------------------

#2;
word <= 'b0111001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1921
#2;

verify(ir === 'b0111, "Assert 7680 : < ir !== 'b0111 >");	// Vector No: 1920
verify(op === 'b11111111, "Assert 7681 : < op !== 'b11111111 >");
verify(extop === 1, "Assert 7682 : < extop !== 1 >");
verify(addr === 'b11111111111111111111, "Assert 7683 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111001111111111111111111111111111111111111111111111111111111111:0:1:1111:11111111:0:11111111111111111111:
//------------------------

#2;
word <= 'b0111001111111111111111111111111111111111111111111111111111111111;
pe <= 0;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1922
#2;

verify(ir === 'b1111, "Assert 7684 : < ir !== 'b1111 >");	// Vector No: 1921
verify(op === 'b11111111, "Assert 7685 : < op !== 'b11111111 >");
verify(extop === 0, "Assert 7686 : < extop !== 0 >");
verify(addr === 'b11111111111111111111, "Assert 7687 : < addr !== 'b11111111111111111111 >");
#2;
clk <= 0;

// 0111001111111111111111111111111111111111111111111111111111111111:1:0:0011:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b0111001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 0;
#2;
clk <= 1;		// Cycle No: 1923
#2;

verify(ir === 'b0011, "Assert 7688 : < ir !== 'b0011 >");	// Vector No: 1922
verify(op === 'b11111000, "Assert 7689 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7690 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7691 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

// 0111001111111111111111111111111111111111111111111111111111111111:1:1:1111:11111000:0:00000111111111111111:
//------------------------

#2;
word <= 'b0111001111111111111111111111111111111111111111111111111111111111;
pe <= 1;
tkk <= 1;
#2;
clk <= 1;		// Cycle No: 1924
#2;

verify(ir === 'b1111, "Assert 7692 : < ir !== 'b1111 >");	// Vector No: 1923
verify(op === 'b11111000, "Assert 7693 : < op !== 'b11111000 >");
verify(extop === 0, "Assert 7694 : < extop !== 0 >");
verify(addr === 'b00000111111111111111, "Assert 7695 : < addr !== 'b00000111111111111111 >");
#2;
clk <= 0;

#4;
if (fail) begin
    $display("Test FAIL");
    $display("------------------------");
    $finish(1);
end
$display("Test PASS");
$display("------------------------");
$finish;

end

endmodule
