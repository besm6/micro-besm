module testbench();

//TODO

endmodule
